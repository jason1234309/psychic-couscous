module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_SING_X0Y150_IOB_X0Y150_IPAD,
  input LIOB33_SING_X0Y199_IOB_X0Y199_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y151_IOB_X0Y151_IPAD,
  input LIOB33_X0Y151_IOB_X0Y152_IPAD,
  input LIOB33_X0Y153_IOB_X0Y153_IPAD,
  input LIOB33_X0Y153_IOB_X0Y154_IPAD,
  input LIOB33_X0Y155_IOB_X0Y155_IPAD,
  input LIOB33_X0Y155_IOB_X0Y156_IPAD,
  input LIOB33_X0Y157_IOB_X0Y157_IPAD,
  input LIOB33_X0Y157_IOB_X0Y158_IPAD,
  input LIOB33_X0Y159_IOB_X0Y159_IPAD,
  input LIOB33_X0Y159_IOB_X0Y160_IPAD,
  input LIOB33_X0Y161_IOB_X0Y161_IPAD,
  input LIOB33_X0Y161_IOB_X0Y162_IPAD,
  input LIOB33_X0Y163_IOB_X0Y163_IPAD,
  input LIOB33_X0Y163_IOB_X0Y164_IPAD,
  input LIOB33_X0Y165_IOB_X0Y165_IPAD,
  input LIOB33_X0Y165_IOB_X0Y166_IPAD,
  input LIOB33_X0Y167_IOB_X0Y167_IPAD,
  input LIOB33_X0Y167_IOB_X0Y168_IPAD,
  input LIOB33_X0Y169_IOB_X0Y169_IPAD,
  input LIOB33_X0Y169_IOB_X0Y170_IPAD,
  input LIOB33_X0Y171_IOB_X0Y171_IPAD,
  input LIOB33_X0Y171_IOB_X0Y172_IPAD,
  input LIOB33_X0Y173_IOB_X0Y173_IPAD,
  input LIOB33_X0Y173_IOB_X0Y174_IPAD,
  input LIOB33_X0Y175_IOB_X0Y175_IPAD,
  input LIOB33_X0Y175_IOB_X0Y176_IPAD,
  input LIOB33_X0Y177_IOB_X0Y177_IPAD,
  input LIOB33_X0Y177_IOB_X0Y178_IPAD,
  input LIOB33_X0Y179_IOB_X0Y179_IPAD,
  input LIOB33_X0Y179_IOB_X0Y180_IPAD,
  input LIOB33_X0Y181_IOB_X0Y181_IPAD,
  input LIOB33_X0Y181_IOB_X0Y182_IPAD,
  input LIOB33_X0Y183_IOB_X0Y183_IPAD,
  input LIOB33_X0Y183_IOB_X0Y184_IPAD,
  input LIOB33_X0Y185_IOB_X0Y185_IPAD,
  input LIOB33_X0Y185_IOB_X0Y186_IPAD,
  input LIOB33_X0Y187_IOB_X0Y187_IPAD,
  input LIOB33_X0Y187_IOB_X0Y188_IPAD,
  input LIOB33_X0Y189_IOB_X0Y189_IPAD,
  input LIOB33_X0Y189_IOB_X0Y190_IPAD,
  input LIOB33_X0Y191_IOB_X0Y191_IPAD,
  input LIOB33_X0Y191_IOB_X0Y192_IPAD,
  input LIOB33_X0Y193_IOB_X0Y193_IPAD,
  input LIOB33_X0Y193_IOB_X0Y194_IPAD,
  input LIOB33_X0Y195_IOB_X0Y195_IPAD,
  input LIOB33_X0Y195_IOB_X0Y196_IPAD,
  input LIOB33_X0Y197_IOB_X0Y197_IPAD,
  input LIOB33_X0Y197_IOB_X0Y198_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y50_IOB_X0Y50_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y51_IOB_X0Y51_OPAD,
  output LIOB33_X0Y51_IOB_X0Y52_OPAD,
  output LIOB33_X0Y53_IOB_X0Y53_OPAD,
  output LIOB33_X0Y53_IOB_X0Y54_OPAD,
  output LIOB33_X0Y55_IOB_X0Y55_OPAD,
  output LIOB33_X0Y55_IOB_X0Y56_OPAD,
  output LIOB33_X0Y57_IOB_X0Y57_OPAD,
  output LIOB33_X0Y57_IOB_X0Y58_OPAD,
  output LIOB33_X0Y59_IOB_X0Y59_OPAD,
  output LIOB33_X0Y59_IOB_X0Y60_OPAD,
  output LIOB33_X0Y61_IOB_X0Y61_OPAD,
  output LIOB33_X0Y61_IOB_X0Y62_OPAD,
  output LIOB33_X0Y63_IOB_X0Y63_OPAD,
  output RIOB33_SING_X105Y149_IOB_X1Y149_OPAD,
  output RIOB33_X105Y123_IOB_X1Y124_OPAD,
  output RIOB33_X105Y125_IOB_X1Y125_OPAD,
  output RIOB33_X105Y125_IOB_X1Y126_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD,
  output RIOB33_X105Y135_IOB_X1Y136_OPAD,
  output RIOB33_X105Y137_IOB_X1Y137_OPAD,
  output RIOB33_X105Y137_IOB_X1Y138_OPAD,
  output RIOB33_X105Y139_IOB_X1Y139_OPAD,
  output RIOB33_X105Y139_IOB_X1Y140_OPAD,
  output RIOB33_X105Y141_IOB_X1Y141_OPAD,
  output RIOB33_X105Y141_IOB_X1Y142_OPAD,
  output RIOB33_X105Y143_IOB_X1Y143_OPAD,
  output RIOB33_X105Y143_IOB_X1Y144_OPAD,
  output RIOB33_X105Y145_IOB_X1Y145_OPAD,
  output RIOB33_X105Y145_IOB_X1Y146_OPAD,
  output RIOB33_X105Y147_IOB_X1Y147_OPAD,
  output RIOB33_X105Y147_IOB_X1Y148_OPAD
  );
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_A;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_A1;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_A2;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_A3;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_A4;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_A5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_A6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_AMUX;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_AO5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_AO6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_A_CY;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_A_XOR;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_B;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_B1;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_B2;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_B3;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_B4;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_B5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_B6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_BMUX;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_BO5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_BO6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_B_CY;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_B_XOR;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_C;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_C1;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_C2;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_C3;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_C4;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_C5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_C6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_CMUX;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_CO5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_CO6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_C_CY;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_C_XOR;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_D;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_D1;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_D2;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_D3;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_D4;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_D5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_D6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_DMUX;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_DO5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_DO6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_D_CY;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X38Y133_D_XOR;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_A;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_A1;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_A2;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_A3;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_A4;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_A5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_A6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_AO5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_AO6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_A_CY;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_A_XOR;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_B;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_B1;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_B2;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_B3;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_B4;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_B5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_B6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_BO5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_BO6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_B_CY;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_B_XOR;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_C;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_C1;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_C2;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_C3;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_C4;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_C5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_C6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_CO5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_CO6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_C_CY;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_C_XOR;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_D;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_D1;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_D2;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_D3;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_D4;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_D5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_D6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_DO5;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_DO6;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_D_CY;
  wire [0:0] CLBLL_L_X26Y133_SLICE_X39Y133_D_XOR;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_A;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_A1;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_A2;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_A3;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_A4;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_A5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_A6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_AMUX;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_AO5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_AO6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_A_CY;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_A_XOR;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_B;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_B1;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_B2;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_B3;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_B4;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_B5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_B6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_BO5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_BO6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_B_CY;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_B_XOR;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_C;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_C1;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_C2;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_C3;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_C4;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_C5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_C6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_CO5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_CO6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_C_CY;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_C_XOR;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_D;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_D1;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_D2;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_D3;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_D4;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_D5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_D6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_DO5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_DO6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_D_CY;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X38Y135_D_XOR;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_A;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_A1;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_A2;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_A3;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_A4;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_A5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_A6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_AO5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_AO6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_A_CY;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_A_XOR;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_B;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_B1;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_B2;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_B3;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_B4;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_B5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_B6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_BO5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_BO6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_B_CY;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_B_XOR;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_C;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_C1;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_C2;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_C3;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_C4;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_C5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_C6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_CO5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_CO6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_C_CY;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_C_XOR;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_D;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_D1;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_D2;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_D3;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_D4;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_D5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_D6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_DO5;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_DO6;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_D_CY;
  wire [0:0] CLBLL_L_X26Y135_SLICE_X39Y135_D_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_AMUX;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_BMUX;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_BO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_BO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_CO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_CO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_DO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_DO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_AO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_AO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_BO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_BO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_CO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_CO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_DO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_DO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D_XOR;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_A;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_A1;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_A2;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_A3;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_A4;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_A5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_A6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_AMUX;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_AO5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_AO6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_A_CY;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_A_XOR;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_B;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_B1;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_B2;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_B3;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_B4;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_B5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_B6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_BO5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_BO6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_B_CY;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_B_XOR;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_C;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_C1;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_C2;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_C3;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_C4;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_C5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_C6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_CO5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_CO6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_C_CY;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_C_XOR;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_D;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_D1;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_D2;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_D3;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_D4;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_D5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_D6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_DO5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_DO6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_D_CY;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X38Y138_D_XOR;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_A;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_A1;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_A2;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_A3;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_A4;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_A5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_A6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_AO5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_AO6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_A_CY;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_A_XOR;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_B;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_B1;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_B2;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_B3;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_B4;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_B5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_B6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_BO5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_BO6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_B_CY;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_B_XOR;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_C;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_C1;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_C2;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_C3;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_C4;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_C5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_C6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_CO5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_CO6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_C_CY;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_C_XOR;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_D;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_D1;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_D2;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_D3;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_D4;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_D5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_D6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_DO5;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_DO6;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_D_CY;
  wire [0:0] CLBLL_L_X26Y138_SLICE_X39Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CLK;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X0Y116_SR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_A_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_B_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_C_XOR;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D1;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D2;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D3;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D4;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO5;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_CY;
  wire [0:0] CLBLL_L_X2Y116_SLICE_X1Y116_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AMUX;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AQ;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AX;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BQ;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BX;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CE;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CLK;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_SR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AQ;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AX;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CE;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CLK;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_SR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_AO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_BO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_BO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_CO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_CO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_DO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_DO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AQ;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AX;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_BO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_BO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CE;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CLK;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_DO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_DO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_SR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AQ;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AX;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CE;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CLK;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_SR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_AO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_AO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_A_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_BO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_BO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_B_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_CO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_CO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_C_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_DO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_DO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X0Y135_D_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A5Q;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_AMUX;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_AO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_AO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_A_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_BO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_BO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_B_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CE;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CLK;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_CO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_C_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D1;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D2;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D3;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D4;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_DO5;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_DO6;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D_CY;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_D_XOR;
  wire [0:0] CLBLL_L_X2Y135_SLICE_X1Y135_SR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_AMUX;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_AO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_AQ;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_AX;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_A_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_BO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_BQ;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_BX;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_B_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_CE;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_CLK;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_CO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_CO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_C_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_DO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_DO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_D_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X0Y137_SR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_AMUX;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_AO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_AO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_A_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_BMUX;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_BO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_BO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_B_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_CO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_CO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_C_XOR;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D1;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D2;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D3;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D4;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_DO5;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_DO6;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D_CY;
  wire [0:0] CLBLL_L_X2Y137_SLICE_X1Y137_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AMUX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BMUX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CMUX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_COUT;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DMUX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AMUX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AQ;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BQ;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CE;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CLK;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_SR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CIN;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_COUT;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_DMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_DO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_DO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_DX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CE;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CLK;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DQ;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_SR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AMUX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AQ;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BMUX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BQ;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CE;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CIN;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CLK;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CMUX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_COUT;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CQ;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_DMUX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_DO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_DO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_DX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_SR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_AO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_AQ;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_AX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_BO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_BO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_BQ;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_BX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CE;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CLK;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_COUT;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CQ;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_DO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_DO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_DQ;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_DX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_SR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AMUX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BMUX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CE;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CIN;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CLK;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CMUX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_COUT;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_DO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_DO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_DX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_SR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AQ;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BQ;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CE;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CIN;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CLK;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_COUT;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CQ;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DMUX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_SR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AX;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_BO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_BO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CE;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CLK;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_DO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_DO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_SR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AQ;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AX;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BQ;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BX;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CE;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CIN;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CLK;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CMUX;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_COUT;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CX;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DMUX;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DX;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_SR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_AO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_AO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_AQ;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_BO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_BO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_CE;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_CLK;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_CO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_CO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_DO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_DO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_SR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_AO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_AO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_AQ;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_AX;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_BO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_BO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_BQ;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_BX;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CE;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CIN;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CLK;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_COUT;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CX;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_DO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_DO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_DX;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_SR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A5Q;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AMUX;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AQ;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_BO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_BO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_BQ;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_BX;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_CE;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_CLK;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_CO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_CO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_DO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_DO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_SR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_AMUX;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_AO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_AO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_BO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_BO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_CO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_CO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_DO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_DO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A5Q;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AMUX;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CE;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CLK;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_SR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CLK;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_SR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A5Q;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AMUX;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AQ;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CE;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CLK;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_SR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AMUX;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CLK;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_SR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_BO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_CO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_DO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_DO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_DO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_DO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AX;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_BO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_BO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CLK;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_DO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_DO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_SR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_CO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_CO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_DO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_DO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A5Q;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AMUX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AQ;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B5Q;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BMUX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BQ;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C5Q;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CE;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CLK;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CMUX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CQ;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D5Q;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DMUX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DQ;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_SR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AMUX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BQ;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CE;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CLK;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_DO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_SR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AQ;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BQ;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CE;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CLK;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_SR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AQ;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CE;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CLK;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_DO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_SR;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_A;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_A1;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_A2;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_A3;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_A4;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_A5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_A6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_AO5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_AO6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_AQ;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_AX;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_A_CY;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_A_XOR;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_B;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_B1;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_B2;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_B3;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_B4;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_B5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_B6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_BO5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_BO6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_BQ;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_BX;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_B_CY;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_B_XOR;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_C;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_C1;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_C2;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_C3;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_C4;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_C5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_C6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_CE;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_CLK;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_CO5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_CO6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_CQ;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_CX;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_C_CY;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_C_XOR;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_D;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_D1;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_D2;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_D3;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_D4;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_D5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_D6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_DO5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_DO6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_DQ;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_DX;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_D_CY;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_D_XOR;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X0Y156_SR;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_A;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_A1;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_A2;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_A3;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_A4;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_A5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_A6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_AO5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_AO6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_A_CY;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_A_XOR;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_B;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_B1;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_B2;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_B3;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_B4;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_B5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_B6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_BO5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_BO6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_B_CY;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_B_XOR;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_C;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_C1;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_C2;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_C3;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_C4;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_C5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_C6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_CO5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_CO6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_C_CY;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_C_XOR;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_D;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_D1;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_D2;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_D3;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_D4;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_D5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_D6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_DO5;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_DO6;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_D_CY;
  wire [0:0] CLBLL_L_X2Y156_SLICE_X1Y156_D_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_AO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_AO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_AQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_AX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_A_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_BMUX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_BO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_BO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_BQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_BX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_B_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CE;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CLK;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_CX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_C_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_DO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_DO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_DQ;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_DX;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_D_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X0Y157_SR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_AO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_AO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_A_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_BO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_BO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_B_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_CO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_CO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_C_XOR;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D1;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D2;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D3;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D4;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_DO5;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_DO6;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D_CY;
  wire [0:0] CLBLL_L_X2Y157_SLICE_X1Y157_D_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A5Q;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_AMUX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_AO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_AO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_AQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_AX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_A_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_BO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_BO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_BQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_BX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_B_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CE;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CLK;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_CX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_C_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_DO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_DO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_DQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_DX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_D_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X0Y158_SR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_AO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_AO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_AQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_AX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_A_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_BO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_BO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_BQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_BX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_B_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_CE;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_CLK;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_CO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_CO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_CQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_CX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_C_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D1;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D2;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D3;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D4;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_DO5;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_DO6;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_DQ;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_DX;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D_CY;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_D_XOR;
  wire [0:0] CLBLL_L_X2Y158_SLICE_X1Y158_SR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CE;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CLK;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_SR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_SR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CE;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_SR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CLK;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_SR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CE;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CLK;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_SR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CE;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CLK;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_SR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CE;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CLK;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_SR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CE;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CLK;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_SR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CLK;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_SR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CLK;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_SR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CLK;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_SR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CLK;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_COUT;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_SR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_F7AMUX_O;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CIN;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_COUT;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_SR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CIN;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_COUT;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_SR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CIN;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CLK;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_COUT;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_SR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CE;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_SR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CE;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_SR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CE;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CLK;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_SR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CE;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CLK;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_SR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CLK;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_SR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CE;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CLK;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_SR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_BO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_BO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_CO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_DO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_DO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CE;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CLK;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_SR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_AO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_AO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_BO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_BO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_DO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_DO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BMUX;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DMUX;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CE;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_SR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_SR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_SR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AMUX;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CLK;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_SR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_SR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CE;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CLK;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_SR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CLK;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_SR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CE;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CLK;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_SR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CE;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CLK;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_SR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CLK;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_SR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CE;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CLK;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_SR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CLK;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_SR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_SR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_SR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_COUT;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CIN;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_COUT;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_SR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CIN;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_COUT;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CIN;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_COUT;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AMUX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BMUX;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CE;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CLK;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X16Y128_SR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_A_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_B_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CLK;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_C_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D1;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D2;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D3;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D4;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO5;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_CY;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_D_XOR;
  wire [0:0] CLBLM_L_X12Y128_SLICE_X17Y128_SR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CLK;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X16Y129_SR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AMUX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_AX;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_A_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_B_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CE;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CLK;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_C_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D1;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D2;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D3;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D4;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO5;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_CY;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_D_XOR;
  wire [0:0] CLBLM_L_X12Y129_SLICE_X17Y129_SR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CE;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X16Y130_SR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AMUX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_AX;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_A_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_B_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CE;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CLK;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_C_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D1;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D2;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D3;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D4;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO5;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_CY;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_D_XOR;
  wire [0:0] CLBLM_L_X12Y130_SLICE_X17Y130_SR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A5Q;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CE;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CLK;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_SR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A5Q;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AMUX;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CE;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CLK;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_SR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A5Q;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B5Q;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CE;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CLK;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_SR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B5Q;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BMUX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CLK;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DMUX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_SR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BMUX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CE;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CLK;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_SR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CLK;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_SR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CLK;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_SR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AX;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CE;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CLK;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_SR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CE;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CLK;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_DO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_SR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CLK;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_DO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_SR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BQ;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CLK;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_SR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BQ;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CLK;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_SR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BI;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CE;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CLK;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_DI;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AQ;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BQ;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CE;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CLK;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_SR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AI;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BI;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CE;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CI;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CLK;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DI;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DMUX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AI;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BI;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CE;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CI;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CLK;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CMUX;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DI;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CLK;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_DMUX;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_DO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_SR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AI;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BI;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CE;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CI;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CLK;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CMUX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_DI;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AMUX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CLK;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_DO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_SR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AI;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BI;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CE;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CI;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CLK;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_DI;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AMUX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CLK;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DMUX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_SR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BMUX;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CLK;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_SR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_F7AMUX_O;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CLK;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_SR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AMUX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CMUX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_F7AMUX_O;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CLK;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_COUT;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_SR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CLK;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_COUT;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_SR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CIN;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_COUT;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CIN;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CLK;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_COUT;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_SR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CIN;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_COUT;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CIN;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CLK;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_COUT;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_SR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AMUX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AMUX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BMUX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CIN;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CLK;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CMUX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_COUT;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_SR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_F7AMUX_O;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_F7BMUX_O;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_A;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_A1;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_A2;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_A3;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_A4;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_A5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_A6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_AO5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_AO6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_AQ;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_A_CY;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_A_XOR;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_B;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_B1;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_B2;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_B3;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_B4;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_B5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_B6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_BO5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_BO6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_B_CY;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_B_XOR;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_C;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_C1;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_C2;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_C3;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_C4;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_C5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_C6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_CE;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_CLK;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_CO5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_CO6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_C_CY;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_C_XOR;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_D;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_D1;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_D2;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_D3;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_D4;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_D5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_D6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_DO5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_DO6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_D_CY;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_D_XOR;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X22Y131_SR;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_A;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_A1;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_A2;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_A3;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_A4;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_A5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_A6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_AO5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_AO6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_A_CY;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_A_XOR;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_B;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_B1;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_B2;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_B3;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_B4;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_B5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_B6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_BO5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_BO6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_B_CY;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_B_XOR;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_C;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_C1;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_C2;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_C3;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_C4;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_C5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_C6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_CO5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_CO6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_C_CY;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_C_XOR;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_D;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_D1;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_D2;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_D3;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_D4;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_D5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_D6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_DO5;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_DO6;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_D_CY;
  wire [0:0] CLBLM_L_X16Y131_SLICE_X23Y131_D_XOR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_A;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_A1;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_A2;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_A3;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_A4;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_A5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_A6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_AO5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_AO6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_AQ;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_A_CY;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_A_XOR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_B;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_B1;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_B2;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_B3;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_B4;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_B5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_B6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_BO5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_BO6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_BQ;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_B_CY;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_B_XOR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_C;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_C1;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_C2;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_C3;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_C4;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_C5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_C6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_CLK;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_CO5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_CO6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_CQ;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_C_CY;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_C_XOR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_D;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_D1;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_D2;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_D3;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_D4;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_D5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_D6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_DO5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_DO6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_D_CY;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_D_XOR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X22Y133_SR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_A;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_A1;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_A2;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_A3;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_A4;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_A5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_A6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_AO5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_AO6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_AQ;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_A_CY;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_A_XOR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_B;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_B1;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_B2;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_B3;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_B4;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_B5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_B6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_BO5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_BO6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_BQ;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_B_CY;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_B_XOR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_C;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_C1;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_C2;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_C3;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_C4;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_C5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_C6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_CLK;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_CO5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_CO6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_CQ;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_C_CY;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_C_XOR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_D;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_D1;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_D2;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_D3;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_D4;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_D5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_D6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_DO5;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_DO6;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_DQ;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_D_CY;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_D_XOR;
  wire [0:0] CLBLM_L_X16Y133_SLICE_X23Y133_SR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_A;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_A1;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_A2;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_A3;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_A4;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_A5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_A6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_AMUX;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_AO5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_AO6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_A_CY;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_A_XOR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_B;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_B1;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_B2;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_B3;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_B4;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_B5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_B6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_BO5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_BO6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_BQ;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_B_CY;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_B_XOR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_C;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_C1;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_C2;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_C3;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_C4;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_C5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_C6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_CLK;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_CO5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_CO6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_C_CY;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_C_XOR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_D;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_D1;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_D2;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_D3;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_D4;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_D5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_D6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_DO5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_DO6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_D_CY;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_D_XOR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X22Y134_SR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_A;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_A1;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_A2;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_A3;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_A4;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_A5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_A6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_AO5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_AO6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_AQ;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_A_CY;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_A_XOR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_B;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_B1;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_B2;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_B3;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_B4;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_B5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_B6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_BO5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_BO6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_B_CY;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_B_XOR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_C;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_C1;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_C2;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_C3;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_C4;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_C5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_C6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_CLK;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_CO5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_CO6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_C_CY;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_C_XOR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_D;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_D1;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_D2;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_D3;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_D4;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_D5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_D6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_DO5;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_DO6;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_D_CY;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_D_XOR;
  wire [0:0] CLBLM_L_X16Y134_SLICE_X23Y134_SR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_AO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_AO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_A_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_BO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_BO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_B_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_CLK;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_CO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_CO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_C_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_DO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_DO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_D_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X22Y135_SR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_AO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_AO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_AQ;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_A_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_BO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_BO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_B_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_CLK;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_CO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_CO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_C_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D1;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D2;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D3;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D4;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_DO5;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_DO6;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D_CY;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_D_XOR;
  wire [0:0] CLBLM_L_X16Y135_SLICE_X23Y135_SR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_AMUX;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_AO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_A_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_BO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_BO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_BQ;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_B_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_CLK;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_CO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_CO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_C_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_DO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_DO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_D_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X22Y136_SR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_AO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_AO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_AQ;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_A_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_BO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_BO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_BQ;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_B_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_CLK;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_CO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_CO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_CQ;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_C_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D1;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D2;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D3;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D4;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_DO5;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_DO6;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_DQ;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D_CY;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_D_XOR;
  wire [0:0] CLBLM_L_X16Y136_SLICE_X23Y136_SR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_AMUX;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_AO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_AO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_A_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_BMUX;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_BO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_BO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_B_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_CO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_CO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_C_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_DO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_DO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X22Y137_D_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_AMUX;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_AO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_AO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_A_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_BO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_BO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_BQ;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_B_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_CLK;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_CO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_CO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_CQ;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_C_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D1;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D2;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D3;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D4;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_DO5;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_DO6;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D_CY;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_D_XOR;
  wire [0:0] CLBLM_L_X16Y137_SLICE_X23Y137_SR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_A;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_A1;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_A2;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_A3;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_A4;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_A5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_A6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_AO5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_AO6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_AQ;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_A_CY;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_A_XOR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_B;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_B1;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_B2;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_B3;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_B4;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_B5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_B6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_BO5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_BO6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_B_CY;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_B_XOR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_C;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_C1;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_C2;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_C3;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_C4;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_C5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_C6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_CLK;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_CO5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_CO6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_C_CY;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_C_XOR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_D;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_D1;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_D2;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_D3;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_D4;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_D5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_D6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_DO5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_DO6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_D_CY;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_D_XOR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X22Y138_SR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_A;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_A1;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_A2;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_A3;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_A4;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_A5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_A6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_AO5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_AO6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_AQ;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_A_CY;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_A_XOR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_B;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_B1;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_B2;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_B3;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_B4;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_B5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_B6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_BO5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_BO6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_B_CY;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_B_XOR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_C;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_C1;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_C2;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_C3;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_C4;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_C5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_C6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_CLK;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_CO5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_CO6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_C_CY;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_C_XOR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_D;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_D1;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_D2;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_D3;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_D4;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_D5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_D6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_DO5;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_DO6;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_D_CY;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_D_XOR;
  wire [0:0] CLBLM_L_X16Y138_SLICE_X23Y138_SR;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_A;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_A1;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_A2;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_A3;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_A4;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_A5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_A6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_AO5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_AO6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_AQ;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_A_CY;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_A_XOR;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_B;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_B1;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_B2;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_B3;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_B4;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_B5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_B6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_BO5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_BO6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_BQ;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_B_CY;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_B_XOR;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_C;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_C1;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_C2;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_C3;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_C4;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_C5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_C6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_CLK;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_CO5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_CO6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_C_CY;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_C_XOR;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_D;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_D1;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_D2;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_D3;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_D4;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_D5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_D6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_DO5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_DO6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_D_CY;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_D_XOR;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X22Y139_SR;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_A;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_A1;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_A2;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_A3;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_A4;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_A5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_A6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_AO5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_AO6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_A_CY;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_A_XOR;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_B;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_B1;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_B2;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_B3;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_B4;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_B5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_B6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_BO5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_BO6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_B_CY;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_B_XOR;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_C;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_C1;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_C2;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_C3;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_C4;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_C5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_C6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_CO5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_CO6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_C_CY;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_C_XOR;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_D;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_D1;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_D2;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_D3;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_D4;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_D5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_D6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_DO5;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_DO6;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_D_CY;
  wire [0:0] CLBLM_L_X16Y139_SLICE_X23Y139_D_XOR;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_A;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_A1;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_A2;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_A3;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_A4;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_A5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_A6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_AO5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_AO6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_AQ;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_AX;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_A_CY;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_A_XOR;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_B;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_B1;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_B2;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_B3;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_B4;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_B5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_B6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_BO5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_BO6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_BQ;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_BX;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_B_CY;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_B_XOR;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_C;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_C1;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_C2;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_C3;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_C4;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_C5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_C6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_CE;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_CLK;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_CO5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_CO6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_CQ;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_CX;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_C_CY;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_C_XOR;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_D;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_D1;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_D2;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_D3;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_D4;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_D5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_D6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_DO5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_DO6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_D_CY;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_D_XOR;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X22Y140_SR;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_A;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_A1;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_A2;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_A3;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_A4;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_A5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_A6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_AO5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_AO6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_A_CY;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_A_XOR;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_B;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_B1;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_B2;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_B3;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_B4;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_B5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_B6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_BO5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_BO6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_B_CY;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_B_XOR;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_C;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_C1;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_C2;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_C3;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_C4;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_C5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_C6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_CO5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_CO6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_C_CY;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_C_XOR;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_D;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_D1;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_D2;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_D3;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_D4;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_D5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_D6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_DO5;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_DO6;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_D_CY;
  wire [0:0] CLBLM_L_X16Y140_SLICE_X23Y140_D_XOR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_A;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_A1;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_A2;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_A3;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_A4;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_A5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_A6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_AMUX;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_AO5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_AO6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_AQ;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_AX;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_A_CY;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_A_XOR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_B;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_B1;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_B2;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_B3;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_B4;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_B5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_B6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_BMUX;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_BO5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_BO6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_BQ;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_BX;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_B_CY;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_B_XOR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_C;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_C1;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_C2;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_C3;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_C4;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_C5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_C6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_CE;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_CLK;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_CO5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_CO6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_CQ;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_CX;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_C_CY;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_C_XOR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_D;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_D1;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_D2;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_D3;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_D4;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_D5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_D6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_DO5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_DO6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_D_CY;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_D_XOR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X22Y141_SR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_A;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_A1;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_A2;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_A3;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_A4;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_A5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_A6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_AO5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_AO6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_AQ;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_AX;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_A_CY;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_A_XOR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_B;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_B1;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_B2;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_B3;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_B4;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_B5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_B6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_BO5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_BO6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_BQ;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_BX;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_B_CY;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_B_XOR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_C;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_C1;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_C2;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_C3;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_C4;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_C5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_C6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_CE;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_CLK;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_CO5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_CO6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_CQ;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_CX;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_C_CY;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_C_XOR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_D;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_D1;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_D2;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_D3;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_D4;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_D5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_D6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_DO5;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_DO6;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_DQ;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_DX;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_D_CY;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_D_XOR;
  wire [0:0] CLBLM_L_X16Y141_SLICE_X23Y141_SR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_A;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_A1;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_A2;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_A3;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_A4;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_A5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_A6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_AMUX;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_AO5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_AO6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_AQ;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_AX;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_A_CY;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_A_XOR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_B;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_B1;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_B2;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_B3;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_B4;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_B5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_B6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_BO5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_BO6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_BQ;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_BX;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_B_CY;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_B_XOR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_C;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_C1;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_C2;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_C3;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_C4;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_C5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_C6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_CE;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_CLK;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_CO5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_CO6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_CQ;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_CX;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_C_CY;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_C_XOR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_D;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_D1;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_D2;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_D3;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_D4;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_D5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_D6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_DO5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_DO6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_DQ;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_DX;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_D_CY;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_D_XOR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X22Y142_SR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_A;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_A1;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_A2;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_A3;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_A4;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_A5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_A6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_AO5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_AO6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_AQ;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_AX;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_A_CY;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_A_XOR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_B;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_B1;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_B2;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_B3;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_B4;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_B5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_B6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_BO5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_BO6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_B_CY;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_B_XOR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_C;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_C1;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_C2;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_C3;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_C4;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_C5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_C6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_CE;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_CLK;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_CO5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_CO6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_C_CY;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_C_XOR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_D;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_D1;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_D2;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_D3;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_D4;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_D5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_D6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_DO5;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_DO6;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_D_CY;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_D_XOR;
  wire [0:0] CLBLM_L_X16Y142_SLICE_X23Y142_SR;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_A;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_A1;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_A2;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_A3;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_A4;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_A5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_A6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_AMUX;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_AO5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_AO6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_AQ;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_AX;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_A_CY;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_A_XOR;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_B;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_B1;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_B2;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_B3;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_B4;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_B5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_B6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_BO5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_BO6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_BQ;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_BX;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_B_CY;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_B_XOR;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_C;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_C1;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_C2;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_C3;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_C4;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_C5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_C6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_CE;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_CLK;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_CO5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_CO6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_CQ;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_CX;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_C_CY;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_C_XOR;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_D;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_D1;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_D2;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_D3;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_D4;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_D5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_D6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_DO5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_DO6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_D_CY;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_D_XOR;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X22Y143_SR;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_A;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_A1;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_A2;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_A3;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_A4;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_A5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_A6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_AO5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_AO6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_A_CY;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_A_XOR;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_B;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_B1;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_B2;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_B3;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_B4;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_B5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_B6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_BO5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_BO6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_B_CY;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_B_XOR;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_C;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_C1;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_C2;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_C3;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_C4;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_C5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_C6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_CO5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_CO6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_C_CY;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_C_XOR;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_D;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_D1;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_D2;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_D3;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_D4;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_D5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_D6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_DO5;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_DO6;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_D_CY;
  wire [0:0] CLBLM_L_X16Y143_SLICE_X23Y143_D_XOR;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_A;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_A1;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_A2;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_A3;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_A4;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_A5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_A6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_AMUX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_AO5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_AO6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_AX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_A_CY;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_A_XOR;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_B;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_B1;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_B2;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_B3;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_B4;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_B5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_B6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_BMUX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_BO5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_BO6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_BX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_B_CY;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_B_XOR;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_C;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_C1;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_C2;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_C3;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_C4;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_C5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_C6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_CMUX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_CO5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_CO6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_COUT;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_CX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_C_CY;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_C_XOR;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_D;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_D1;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_D2;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_D3;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_D4;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_D5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_D6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_DMUX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_DO5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_DO6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_DX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_D_CY;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X22Y150_D_XOR;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_A;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_A1;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_A2;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_A3;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_A4;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_A5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_A6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_AMUX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_AO5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_AO6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_A_CY;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_A_XOR;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_B;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_B1;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_B2;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_B3;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_B4;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_B5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_B6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_BMUX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_BO5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_BO6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_B_CY;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_B_XOR;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_C;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_C1;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_C2;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_C3;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_C4;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_C5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_C6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_CMUX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_CO5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_CO6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_C_CY;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_C_XOR;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_D;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_D1;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_D2;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_D3;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_D4;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_D5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_D6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_DMUX;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_DO5;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_DO6;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_D_CY;
  wire [0:0] CLBLM_L_X16Y150_SLICE_X23Y150_D_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_AMUX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_AO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_AO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_AX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_A_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_BMUX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_BO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_BO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_BX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CIN;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CMUX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_COUT;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_CX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_C_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_DMUX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_DO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_DO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_DX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_AO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_AO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_AQ;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_AX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_A_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_BO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_BO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_B_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_CLK;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_CMUX;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_CO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_CO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_C_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D1;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D2;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D3;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D4;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_DO5;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_DO6;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D_CY;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_D_XOR;
  wire [0:0] CLBLM_L_X16Y151_SLICE_X23Y151_SR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AMUX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_A_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BMUX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_BX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_B_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CMUX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_COUT;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_CX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_C_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_DMUX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_DO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_DO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_DX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X22Y152_D_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_AO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_AO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_AQ;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_A_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_BO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_BO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_B_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_CLK;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_CO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_CO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_C_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D1;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D2;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D3;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D4;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_DMUX;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_DO5;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_DO6;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D_CY;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_D_XOR;
  wire [0:0] CLBLM_L_X16Y152_SLICE_X23Y152_SR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_AMUX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_AO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_AO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_AX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_A_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_BMUX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_BO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_BO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_BX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_B_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_CIN;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_CMUX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_CO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_CO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_COUT;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_CX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_C_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_DMUX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_DO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_DO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_DX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X22Y153_D_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_AMUX;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_AO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_A_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_BO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_BO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_B_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_CO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_CO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_C_XOR;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D1;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D2;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D3;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D4;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_DO5;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_DO6;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D_CY;
  wire [0:0] CLBLM_L_X16Y153_SLICE_X23Y153_D_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_AMUX;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_AO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_AO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_AX;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_A_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_BO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_BO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_BX;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_B_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_CIN;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_CO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_CO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_COUT;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_CX;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_C_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_DO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_DO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_DX;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X22Y154_D_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_AO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_AO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_A_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_BO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_BO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_B_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_CO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_CO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_C_XOR;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D1;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D2;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D3;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D4;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_DO5;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_DO6;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D_CY;
  wire [0:0] CLBLM_L_X16Y154_SLICE_X23Y154_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CE;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_SR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_SR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_SR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_SR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_F7AMUX_O;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_F7BMUX_O;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_F8MUX_O;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_SR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_SR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CLK;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_SR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CLK;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_SR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CLK;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_SR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CLK;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_SR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_SR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CE;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_SR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_SR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_SR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5Q;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_SR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_SR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_SR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_SR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CE;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_SR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CE;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_SR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CE;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_SR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_F7AMUX_O;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CE;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_SR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CE;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_SR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_COUT;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_COUT;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CIN;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_COUT;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CIN;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_COUT;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CE;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CIN;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CLK;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_COUT;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_SR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CIN;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_COUT;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CIN;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_COUT;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CIN;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_COUT;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CE;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CLK;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CMUX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_SR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CLK;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_SR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CLK;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_SR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AMUX;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CLK;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_SR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CE;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CLK;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_SR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CLK;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CMUX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_SR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_F7AMUX_O;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_F7BMUX_O;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_F8MUX_O;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BI;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CE;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CLK;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DI;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CLK;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_SR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BI;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CE;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CLK;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DI;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CE;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CLK;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_SR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AI;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BI;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CE;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CI;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CLK;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DI;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CE;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CLK;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_SR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AI;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BI;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CE;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CI;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DI;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_SR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AI;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BI;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CE;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CI;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CLK;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DI;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AMUX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BMUX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CLK;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CMUX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_F7AMUX_O;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_F7BMUX_O;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_F8MUX_O;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_SR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BMUX;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A5Q;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AMUX;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AX;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CLK;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_SR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CLK;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_SR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CLK;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_SR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CLK;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_SR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A5Q;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AMUX;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B5Q;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BMUX;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CE;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CLK;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X18Y128_SR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_A_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_B_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_C_XOR;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D1;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D2;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D3;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D4;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO5;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_CY;
  wire [0:0] CLBLM_R_X13Y128_SLICE_X19Y128_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B5Q;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BMUX;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CE;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CLK;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_CQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X18Y129_SR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_A_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BMUX;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_B_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CLK;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_C_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D1;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D2;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D3;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D4;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO5;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_CY;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_D_XOR;
  wire [0:0] CLBLM_R_X13Y129_SLICE_X19Y129_SR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CE;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CLK;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X18Y130_SR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_A_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_B_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CLK;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_C_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D1;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D2;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D3;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D4;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO5;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_CY;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_D_XOR;
  wire [0:0] CLBLM_R_X13Y130_SLICE_X19Y130_SR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_AX;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_A_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_BX;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_B_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CE;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CLK;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CMUX;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_CX;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_C_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_DX;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_D_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X18Y131_SR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_A_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_BO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_BQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_B_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CE;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CLK;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_CQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_C_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D1;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D2;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D3;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D4;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_DO5;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_DQ;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D_CY;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_D_XOR;
  wire [0:0] CLBLM_R_X13Y131_SLICE_X19Y131_SR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AMUX;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BMUX;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CLK;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CMUX;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D5Q;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DMUX;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_D_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X18Y132_SR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_A_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_B_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_C_XOR;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D1;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D2;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D3;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D4;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO5;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_CY;
  wire [0:0] CLBLM_R_X13Y132_SLICE_X19Y132_D_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_AMUX;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_AO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_BMUX;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_BO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_CO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_CO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_DO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_DO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A5Q;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_AMUX;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_AO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_AO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_AQ;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B5Q;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_BMUX;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_BO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_BO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_BQ;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_CE;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_CLK;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_CMUX;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_DO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_DO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_SR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_BMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_CO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A5Q;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AQ;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B5Q;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CE;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CLK;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_SR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AMUX;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AX;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_BO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_BO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_BX;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_CE;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_CLK;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_CO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_CO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_DO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_DO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_SR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_AO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_AO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_AQ;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_AX;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_BO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_BO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_BQ;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_BX;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CE;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CLK;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CQ;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CX;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_DO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_DO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_DQ;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_DX;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_SR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A5Q;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AMUX;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B5Q;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_BMUX;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_BO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_BO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_BQ;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CE;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CLK;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_DO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_DO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_SR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_AO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_AO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_AQ;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_BO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_BO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_BQ;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_CLK;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_CO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_CO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_DO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_DO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_SR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AX;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_BO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_BO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CE;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CLK;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_DO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_DO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_SR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_AMUX;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_AO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_AO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_BO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_BO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_BQ;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_CLK;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_CO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_CO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_DO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_DO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_SR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A5Q;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AMUX;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AQ;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_BO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_CE;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_CLK;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_CO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_CO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_DO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_DO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_SR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_AO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_AO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_AQ;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_BO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_BO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_BQ;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_CLK;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_CO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_CO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_CQ;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_DO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_SR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_BI;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_CE;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_CLK;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_DI;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_DO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_AMUX;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_BO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_CO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_CO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_DO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_AI;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_AO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_BI;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_BMUX;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_BO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CE;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CI;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CLK;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_DI;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_DO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_AMUX;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_BMUX;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_BO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_BO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_CO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_CO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_DO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_DO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_BMUX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_CO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_DO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_DO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_BO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_BO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_BQ;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_BX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CE;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CLK;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CQ;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_DO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_DO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_SR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_AO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_BO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_BO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_CO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_CO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_DO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_DO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_AO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_AO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_BO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_BO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_CO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_CO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_DO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_DO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_AMUX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_AO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_AX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_BMUX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_BO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_BO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_BX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_CMUX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_CO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_COUT;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_CX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_DMUX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_DO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_DO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_DX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_AMUX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_AO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_AO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_AX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_BO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_BO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_CMUX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_CO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_CO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_DO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_DO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_AMUX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_AO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_AO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_AX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_BMUX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_BO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_BO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_BX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CIN;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CMUX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_COUT;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_DMUX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_DO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_DO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_DX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_AMUX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_AO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_AO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_BMUX;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_BO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_BO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_CO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_DO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AMUX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_AX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_A_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_BMUX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_BO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_BX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_B_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CIN;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CMUX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_COUT;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_CX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_C_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_DMUX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_DO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_DX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X18Y146_D_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_AMUX;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_AO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_A_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_BO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_BO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_B_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_CO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_CO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_C_XOR;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D1;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D2;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D3;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D4;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_DO5;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_DO6;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D_CY;
  wire [0:0] CLBLM_R_X13Y146_SLICE_X19Y146_D_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AMUX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BMUX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CIN;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CMUX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_COUT;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_DO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_DO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_DX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_AMUX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_AO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_BO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_CMUX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_CO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_CO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_DMUX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_DO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_DO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AMUX;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_BO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_BO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_DO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_AO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_AO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_BO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_BO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_CO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_CO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_DO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_DO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AMUX;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AX;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_DO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_F7AMUX_O;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AMUX;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_BO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_BO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_DO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_DO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_AO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_BO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_CO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_CO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_DO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_DO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_AMUX;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_AO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_AO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_AX;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_BO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_BO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_CO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_CO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_DO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_DO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_F7AMUX_O;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A5Q;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_AMUX;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_AO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_A_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B5Q;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_BMUX;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_BO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_BO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_BQ;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_B_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_CLK;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_CO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_CQ;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_C_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_DO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_D_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X20Y128_SR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_AO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_AO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_A_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_BO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_B_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_CO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_C_XOR;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D1;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D2;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D3;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D4;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_DO5;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_DO6;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D_CY;
  wire [0:0] CLBLM_R_X15Y128_SLICE_X21Y128_D_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_AO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_AO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_AQ;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_A_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_BO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_BO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_BQ;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_B_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CE;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CLK;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_CQ;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_C_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_DO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_DO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_D_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X20Y129_SR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_AO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_AO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_AQ;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_A_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B5Q;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_BMUX;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_BO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_BQ;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_B_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CE;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CLK;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_CQ;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_C_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D1;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D2;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D3;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D4;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_DO5;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D_CY;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_D_XOR;
  wire [0:0] CLBLM_R_X15Y129_SLICE_X21Y129_SR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AMUX;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_AX;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_A_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_BO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_BO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_B_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CE;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CLK;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_CO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_C_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_DO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_DO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_D_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X20Y130_SR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_AO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_AO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_A_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_BO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_BO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_BQ;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_B_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CE;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CLK;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_CQ;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_C_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D1;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D2;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D3;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D4;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_DO5;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_DO6;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D_CY;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_D_XOR;
  wire [0:0] CLBLM_R_X15Y130_SLICE_X21Y130_SR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_AO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_AO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_AQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_A_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_BO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_BO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_BQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_B_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_CE;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_CLK;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_CO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_CO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_CQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_C_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_DO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_DO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_DQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_D_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X20Y131_SR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AMUX;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_AX;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_A_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_BMUX;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_BO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_B_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_CE;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_CLK;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_CO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_CO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_CQ;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_C_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D1;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D2;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D3;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D4;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_DO5;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_DO6;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D_CY;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_D_XOR;
  wire [0:0] CLBLM_R_X15Y131_SLICE_X21Y131_SR;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_A;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_A1;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_A2;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_A3;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_A4;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_A5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_A6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_AO5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_AO6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_A_CY;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_A_XOR;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_B;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_B1;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_B2;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_B3;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_B4;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_B5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_B6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_BO5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_BO6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_B_CY;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_B_XOR;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_C;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_C1;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_C2;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_C3;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_C4;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_C5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_C6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_CO5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_CO6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_C_CY;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_C_XOR;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_D;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_D1;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_D2;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_D3;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_D4;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_D5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_D6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_DO5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_DO6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_D_CY;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X20Y133_D_XOR;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_A;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_A1;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_A2;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_A3;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_A4;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_A5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_A6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_AO5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_AO6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_AQ;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_A_CY;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_A_XOR;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_B;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_B1;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_B2;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_B3;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_B4;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_B5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_B6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_BO5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_BO6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_BQ;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_B_CY;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_B_XOR;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_C;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_C1;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_C2;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_C3;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_C4;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_C5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_C6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_CE;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_CLK;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_CO5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_CO6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_CQ;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_C_CY;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_C_XOR;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_D;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_D1;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_D2;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_D3;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_D4;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_D5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_D6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_DO5;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_DO6;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_D_CY;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_D_XOR;
  wire [0:0] CLBLM_R_X15Y133_SLICE_X21Y133_SR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_A;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_A1;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_A2;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_A3;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_A4;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_A5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_A6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_AMUX;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_AO5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_AO6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_AX;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_A_CY;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_A_XOR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_B;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_B1;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_B2;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_B3;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_B4;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_B5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_B6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_BMUX;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_BO5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_BO6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_BQ;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_BX;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_B_CY;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_B_XOR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_C;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_C1;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_C2;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_C3;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_C4;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_C5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_C6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_CE;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_CLK;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_CMUX;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_CO5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_CO6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_COUT;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_CQ;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_CX;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_C_CY;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_C_XOR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_D;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_D1;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_D2;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_D3;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_D4;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_D5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_D6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_DMUX;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_DO5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_DO6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_DQ;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_DX;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_D_CY;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_D_XOR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X20Y134_SR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_A;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_A1;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_A2;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_A3;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_A4;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_A5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_A6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_AO5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_AO6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_AQ;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_A_CY;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_A_XOR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_B;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_B1;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_B2;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_B3;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_B4;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_B5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_B6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_BO5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_BO6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_BQ;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_B_CY;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_B_XOR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_C;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_C1;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_C2;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_C3;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_C4;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_C5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_C6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_CE;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_CLK;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_CO5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_CO6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_CQ;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_C_CY;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_C_XOR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_D;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_D1;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_D2;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_D3;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_D4;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_D5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_D6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_DO5;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_DO6;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_D_CY;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_D_XOR;
  wire [0:0] CLBLM_R_X15Y134_SLICE_X21Y134_SR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_AMUX;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_AO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_AO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_AX;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_A_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_BMUX;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_BO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_BO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_BX;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_B_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_CIN;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_CMUX;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_CO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_CO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_COUT;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_CX;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_C_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_DMUX;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_DO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_DO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_DX;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X20Y135_D_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_AO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_AO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_AQ;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_A_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_BO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_BO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_BQ;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_B_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_CE;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_CLK;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_CO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_CO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_C_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D1;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D2;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D3;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D4;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_DMUX;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_DO5;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_DO6;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D_CY;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_D_XOR;
  wire [0:0] CLBLM_R_X15Y135_SLICE_X21Y135_SR;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_A;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_A1;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_A2;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_A3;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_A4;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_A5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_A6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_AMUX;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_AO5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_AO6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_AX;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_A_CY;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_A_XOR;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_B;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_B1;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_B2;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_B3;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_B4;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_B5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_B6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_BMUX;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_BO5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_BO6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_BX;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_B_CY;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_B_XOR;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_C;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_C1;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_C2;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_C3;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_C4;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_C5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_C6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_CIN;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_CMUX;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_CO5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_CO6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_COUT;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_CX;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_C_CY;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_C_XOR;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_D;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_D1;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_D2;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_D3;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_D4;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_D5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_D6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_DMUX;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_DO5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_DO6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_DX;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_D_CY;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X20Y136_D_XOR;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_A;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_A1;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_A2;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_A3;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_A4;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_A5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_A6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_AO5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_AO6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_AQ;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_A_CY;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_A_XOR;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_B;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_B1;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_B2;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_B3;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_B4;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_B5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_B6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_BO5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_BO6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_BQ;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_B_CY;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_B_XOR;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_C;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_C1;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_C2;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_C3;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_C4;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_C5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_C6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_CE;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_CLK;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_CO5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_CO6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_CQ;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_C_CY;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_C_XOR;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_D;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_D1;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_D2;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_D3;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_D4;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_D5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_D6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_DO5;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_DO6;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_DQ;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_D_CY;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_D_XOR;
  wire [0:0] CLBLM_R_X15Y136_SLICE_X21Y136_SR;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_A;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_A1;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_A2;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_A3;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_A4;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_A5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_A6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_AMUX;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_AO5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_AO6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_AX;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_A_CY;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_A_XOR;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_B;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_B1;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_B2;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_B3;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_B4;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_B5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_B6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_BMUX;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_BO5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_BO6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_BX;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_B_CY;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_B_XOR;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_C;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_C1;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_C2;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_C3;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_C4;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_C5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_C6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_CIN;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_CMUX;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_CO5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_CO6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_COUT;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_CX;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_C_CY;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_C_XOR;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_D;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_D1;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_D2;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_D3;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_D4;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_D5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_D6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_DMUX;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_DO5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_DO6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_DX;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_D_CY;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X20Y137_D_XOR;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_A;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_A1;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_A2;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_A3;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_A4;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_A5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_A6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_AO5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_AO6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_AQ;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_A_CY;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_A_XOR;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_B;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_B1;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_B2;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_B3;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_B4;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_B5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_B6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_BO5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_BO6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_BQ;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_B_CY;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_B_XOR;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_C;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_C1;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_C2;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_C3;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_C4;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_C5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_C6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_CE;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_CLK;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_CO5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_CO6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_C_CY;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_C_XOR;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_D;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_D1;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_D2;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_D3;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_D4;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_D5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_D6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_DO5;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_DO6;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_D_CY;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_D_XOR;
  wire [0:0] CLBLM_R_X15Y137_SLICE_X21Y137_SR;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_A;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_A1;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_A2;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_A3;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_A4;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_A5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_A6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_AO5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_AO6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_A_CY;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_A_XOR;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_B;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_B1;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_B2;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_B3;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_B4;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_B5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_B6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_BO5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_BO6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_B_CY;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_B_XOR;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_C;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_C1;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_C2;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_C3;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_C4;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_C5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_C6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_CO5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_CO6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_C_CY;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_C_XOR;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_D;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_D1;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_D2;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_D3;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_D4;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_D5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_D6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_DO5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_DO6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_D_CY;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X20Y138_D_XOR;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_A;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_A1;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_A2;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_A3;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_A4;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_A5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_A6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_AO5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_AO6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_AQ;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_A_CY;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_A_XOR;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_B;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_B1;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_B2;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_B3;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_B4;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_B5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_B6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_BO5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_BO6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_BQ;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_B_CY;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_B_XOR;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_C;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_C1;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_C2;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_C3;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_C4;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_C5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_C6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_CE;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_CLK;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_CO5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_CO6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_C_CY;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_C_XOR;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_D;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_D1;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_D2;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_D3;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_D4;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_D5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_D6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_DO5;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_DO6;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_D_CY;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_D_XOR;
  wire [0:0] CLBLM_R_X15Y138_SLICE_X21Y138_SR;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_A;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_A1;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_A2;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_A3;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_A4;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_A5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_A6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_AO5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_AO6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_A_CY;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_A_XOR;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_B;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_B1;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_B2;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_B3;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_B4;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_B5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_B6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_BO5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_BO6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_B_CY;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_B_XOR;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_C;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_C1;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_C2;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_C3;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_C4;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_C5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_C6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_CO5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_CO6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_C_CY;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_C_XOR;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_D;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_D1;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_D2;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_D3;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_D4;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_D5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_D6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_DO5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_DO6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_D_CY;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X20Y139_D_XOR;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_A;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_A1;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_A2;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_A3;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_A4;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_A5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_A6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_AMUX;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_AO5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_AQ;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_AX;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_A_CY;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_A_XOR;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_B;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_B1;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_B2;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_B3;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_B4;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_B5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_B6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_BMUX;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_BO5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_BO6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_BQ;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_BX;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_B_CY;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_B_XOR;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_C;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_C1;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_C2;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_C3;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_C4;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_C5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_C6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_CE;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_CLK;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_CO5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_CO6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_CQ;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_CX;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_C_CY;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_C_XOR;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_D;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_D1;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_D2;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_D3;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_D4;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_D5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_D6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_DO5;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_DO6;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_D_CY;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_D_XOR;
  wire [0:0] CLBLM_R_X15Y139_SLICE_X21Y139_SR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_A;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_A1;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_A2;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_A3;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_A4;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_A5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_A6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_AO5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_AO6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_AQ;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_AX;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_A_CY;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_A_XOR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_B;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_B1;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_B2;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_B3;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_B4;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_B5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_B6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_BO5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_BO6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_BQ;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_BX;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_B_CY;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_B_XOR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_C;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_C1;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_C2;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_C3;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_C4;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_C5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_C6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_CE;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_CLK;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_CO5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_CO6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_CQ;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_CX;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_C_CY;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_C_XOR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_D;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_D1;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_D2;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_D3;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_D4;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_D5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_D6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_DO5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_DO6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_D_CY;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_D_XOR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X20Y140_SR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_A;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_A1;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_A2;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_A3;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_A4;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_A5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_A6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_AMUX;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_AO5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_AQ;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_AX;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_A_CY;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_A_XOR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_B;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_B1;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_B2;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_B3;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_B4;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_B5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_B6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_BO5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_BO6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_BQ;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_BX;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_B_CY;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_B_XOR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_C;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_C1;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_C2;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_C3;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_C4;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_C5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_C6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_CE;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_CLK;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_CMUX;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_CO5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_CO6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_CQ;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_CX;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_C_CY;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_C_XOR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_D;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_D1;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_D2;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_D3;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_D4;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_D5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_D6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_DO5;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_DO6;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_DQ;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_DX;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_D_CY;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_D_XOR;
  wire [0:0] CLBLM_R_X15Y140_SLICE_X21Y140_SR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_A;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_A1;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_A2;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_A3;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_A4;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_A5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_A6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_AO5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_AO6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_AQ;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_AX;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_A_CY;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_A_XOR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_B;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_B1;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_B2;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_B3;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_B4;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_B5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_B6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_BO5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_BO6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_BQ;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_BX;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_B_CY;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_B_XOR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_C;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_C1;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_C2;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_C3;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_C4;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_C5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_C6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_CE;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_CLK;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_CO5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_CO6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_CQ;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_CX;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_C_CY;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_C_XOR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_D;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_D1;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_D2;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_D3;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_D4;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_D5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_D6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_DO5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_DO6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_DQ;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_DX;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_D_CY;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_D_XOR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X20Y141_SR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A1;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A2;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A3;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A4;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A5Q;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_AMUX;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_AO5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_AO6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_AQ;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_AX;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A_CY;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_A_XOR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_B;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_B1;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_B2;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_B3;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_B4;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_B5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_B6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_BO5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_BO6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_BQ;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_BX;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_B_CY;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_B_XOR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_C;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_C1;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_C2;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_C3;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_C4;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_C5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_C6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_CE;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_CLK;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_CO5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_CO6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_CQ;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_CX;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_C_CY;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_C_XOR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_D;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_D1;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_D2;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_D3;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_D4;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_D5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_D6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_DO5;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_DO6;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_DQ;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_DX;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_D_CY;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_D_XOR;
  wire [0:0] CLBLM_R_X15Y141_SLICE_X21Y141_SR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_AMUX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_AO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_AX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_BMUX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_BO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_BO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_BQ;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_BX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C5Q;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CE;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CLK;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CMUX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CQ;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_DO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_DQ;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_DX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_SR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A5Q;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_AMUX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_AO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_AO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_AQ;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_AX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_BO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_BO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_BQ;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_BX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_CE;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_CLK;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_CMUX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_CO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_CO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_CQ;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_CX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_DMUX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_DO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_DO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_DQ;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_DX;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_SR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_A;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_A1;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_A2;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_A3;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_A4;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_A5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_A6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_AMUX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_AO5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_AO6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_AQ;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_AX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_A_CY;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_A_XOR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_B;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_B1;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_B2;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_B3;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_B4;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_B5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_B6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_BO5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_BO6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_BQ;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_BX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_B_CY;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_B_XOR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_C;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_C1;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_C2;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_C3;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_C4;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_C5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_C6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_CE;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_CLK;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_CO5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_CO6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_CQ;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_CX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_C_CY;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_C_XOR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_D;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_D1;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_D2;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_D3;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_D4;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_D5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_D6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_DO5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_DO6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_DQ;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_DX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_D_CY;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_D_XOR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X20Y143_SR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_A;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_A1;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_A2;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_A3;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_A4;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_A5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_A6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_AMUX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_AO6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_AQ;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_AX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_A_CY;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_A_XOR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B1;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B2;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B3;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B4;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B5Q;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_BMUX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_BO5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_BO6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_BQ;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_BX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B_CY;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_B_XOR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_C;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_C1;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_C2;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_C3;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_C4;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_C5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_C6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_CE;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_CLK;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_CMUX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_CO5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_CO6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_CQ;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_CX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_C_CY;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_C_XOR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_D;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_D1;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_D2;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_D3;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_D4;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_D5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_D6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_DO5;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_DO6;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_DQ;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_DX;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_D_CY;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_D_XOR;
  wire [0:0] CLBLM_R_X15Y143_SLICE_X21Y143_SR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_AMUX;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_AO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_AO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_AX;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_A_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_BO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_BO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_BQ;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_BX;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_B_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_CE;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_CLK;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_CO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_CQ;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_CX;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_C_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_DO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_DO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_D_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X20Y144_SR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_AO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_AQ;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_AX;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_A_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_BO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_BQ;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_BX;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_B_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_CE;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_CLK;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_CO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_CQ;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_CX;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_C_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D1;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D2;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D3;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D4;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_DO5;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_DO6;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D_CY;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_D_XOR;
  wire [0:0] CLBLM_R_X15Y144_SLICE_X21Y144_SR;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_A;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_A1;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_A2;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_A3;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_A4;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_A5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_A6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_AMUX;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_AO5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_AO6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_AX;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_A_CY;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_A_XOR;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_B;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_B1;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_B2;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_B3;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_B4;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_B5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_B6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_BO5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_BO6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_B_CY;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_B_XOR;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_C;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_C1;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_C2;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_C3;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_C4;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_C5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_C6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_CO5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_C_CY;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_C_XOR;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_D;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_D1;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_D2;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_D3;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_D4;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_D5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_D6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_DO5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_DO6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_D_CY;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_D_XOR;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_A;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_A1;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_A2;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_A3;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_A4;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_A5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_A6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_AO5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_AO6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_A_CY;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_A_XOR;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_B;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_B1;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_B2;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_B3;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_B4;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_B5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_B6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_BO5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_BO6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_B_CY;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_B_XOR;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_C;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_C1;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_C2;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_C3;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_C4;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_C5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_C6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_CO5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_CO6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_C_CY;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_C_XOR;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_D;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_D1;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_D2;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_D3;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_D4;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_D5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_D6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_DO5;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_DO6;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_D_CY;
  wire [0:0] CLBLM_R_X15Y145_SLICE_X21Y145_D_XOR;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_A;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_A1;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_A2;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_A3;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_A4;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_A5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_A6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_AO5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_A_CY;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_A_XOR;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_B;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_B1;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_B2;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_B3;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_B4;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_B5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_B6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_BO5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_BO6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_B_CY;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_B_XOR;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_C;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_C1;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_C2;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_C3;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_C4;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_C5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_C6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_CO5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_CO6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_C_CY;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_C_XOR;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_D;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_D1;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_D2;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_D3;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_D4;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_D5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_D6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_DO5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_DO6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_D_CY;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X20Y146_D_XOR;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_A;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_A1;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_A2;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_A3;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_A4;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_A5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_A6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_AMUX;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_AO5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_AO6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_AX;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_A_CY;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_A_XOR;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_B;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_B1;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_B2;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_B3;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_B4;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_B5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_B6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_BO5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_BO6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_B_CY;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_B_XOR;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_C;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_C1;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_C2;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_C3;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_C4;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_C5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_C6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_CMUX;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_CO5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_CO6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_C_CY;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_C_XOR;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_D;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_D1;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_D2;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_D3;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_D4;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_D5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_D6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_DO5;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_DO6;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_D_CY;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_D_XOR;
  wire [0:0] CLBLM_R_X15Y146_SLICE_X21Y146_F7AMUX_O;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_A;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_A1;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_A2;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_A3;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_A4;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_A5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_A6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_AO5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_AO6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_A_CY;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_A_XOR;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_B;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_B1;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_B2;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_B3;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_B4;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_B5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_B6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_BO5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_BO6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_B_CY;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_B_XOR;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_C;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_C1;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_C2;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_C3;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_C4;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_C5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_C6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_CO5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_CO6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_C_CY;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_C_XOR;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_D;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_D1;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_D2;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_D3;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_D4;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_D5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_D6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_DO5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_DO6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_D_CY;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X20Y147_D_XOR;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_A;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_A1;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_A2;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_A3;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_A4;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_A5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_A6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_AO5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_AO6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_A_CY;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_A_XOR;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_B;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_B1;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_B2;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_B3;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_B4;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_B5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_B6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_BO5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_BO6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_B_CY;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_B_XOR;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_C;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_C1;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_C2;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_C3;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_C4;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_C5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_C6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_CO5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_CO6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_C_CY;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_C_XOR;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_D;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_D1;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_D2;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_D3;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_D4;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_D5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_D6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_DO5;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_DO6;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_D_CY;
  wire [0:0] CLBLM_R_X15Y147_SLICE_X21Y147_D_XOR;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_A;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_A1;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_A2;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_A3;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_A4;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_A5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_A6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_AO5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_AO6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_A_CY;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_A_XOR;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_B;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_B1;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_B2;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_B3;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_B4;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_B5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_B6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_BMUX;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_BO5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_BO6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_B_CY;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_B_XOR;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_C;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_C1;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_C2;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_C3;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_C4;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_C5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_C6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_CO5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_CO6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_C_CY;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_C_XOR;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_D;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_D1;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_D2;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_D3;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_D4;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_D5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_D6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_DO5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_DO6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_D_CY;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X20Y148_D_XOR;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_A;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_A1;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_A2;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_A3;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_A4;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_A5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_A6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_AMUX;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_AO5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_AO6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_A_CY;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_A_XOR;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_B;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_B1;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_B2;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_B3;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_B4;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_B5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_B6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_BO5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_B_CY;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_B_XOR;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_C;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_C1;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_C2;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_C3;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_C4;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_C5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_C6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_CO5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_CO6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_C_CY;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_C_XOR;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_D;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_D1;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_D2;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_D3;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_D4;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_D5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_D6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_DO5;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_DO6;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_D_CY;
  wire [0:0] CLBLM_R_X15Y148_SLICE_X21Y148_D_XOR;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_A;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_A1;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_A2;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_A3;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_A4;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_A5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_A6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_AMUX;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_AO5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_AO6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_A_CY;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_A_XOR;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_B;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_B1;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_B2;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_B3;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_B4;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_B5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_B6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_BMUX;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_BO5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_BO6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_B_CY;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_B_XOR;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_C;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_C1;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_C2;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_C3;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_C4;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_C5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_C6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_CO5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_CO6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_C_CY;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_C_XOR;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_D;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_D1;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_D2;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_D3;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_D4;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_D5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_D6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_DO5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_DO6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_D_CY;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X20Y149_D_XOR;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_A;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_A1;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_A2;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_A3;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_A4;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_A5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_A6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_AO5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_AO6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_A_CY;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_A_XOR;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_B;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_B1;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_B2;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_B3;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_B4;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_B5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_B6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_BO5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_BO6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_B_CY;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_B_XOR;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_C;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_C1;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_C2;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_C3;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_C4;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_C5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_C6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_CO5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_CO6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_C_CY;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_C_XOR;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_D;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_D1;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_D2;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_D3;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_D4;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_D5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_D6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_DO5;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_DO6;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_D_CY;
  wire [0:0] CLBLM_R_X15Y149_SLICE_X21Y149_D_XOR;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_A;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_A1;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_A2;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_A3;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_A4;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_A5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_A6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_AO5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_AO6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_A_CY;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_A_XOR;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_B;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_B1;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_B2;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_B3;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_B4;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_B5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_B6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_BO5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_BO6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_B_CY;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_B_XOR;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_C;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_C1;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_C2;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_C3;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_C4;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_C5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_C6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_CLK;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_CO5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_CO6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_C_CY;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_C_XOR;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_D;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_D1;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_D2;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_D3;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_D4;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_D5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_D6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_DMUX;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_D_CY;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_D_XOR;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X20Y150_SR;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_A;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_A1;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_A2;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_A3;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_A4;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_A5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_A6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_AMUX;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_AO5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_AO6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_A_CY;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_A_XOR;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_B;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_B1;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_B2;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_B3;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_B4;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_B5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_B6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_BO5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_BO6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_B_CY;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_B_XOR;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_C;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_C1;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_C2;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_C3;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_C4;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_C5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_C6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_CMUX;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_CO5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_CO6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_C_CY;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_C_XOR;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_D;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_D1;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_D2;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_D3;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_D4;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_D5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_D6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_DO5;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_DO6;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_D_CY;
  wire [0:0] CLBLM_R_X15Y150_SLICE_X21Y150_D_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AMUX;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AX;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_BMUX;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_BO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_BO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_BQ;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_BX;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CLK;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CMUX;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_DO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_SR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A5Q;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_AMUX;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_AO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_AO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_AX;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_BMUX;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_BO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_CLK;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_CO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_CO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_DO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_SR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_A;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_A1;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_A2;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_A3;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_A4;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_A5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_A6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_AO5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_AO6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_AQ;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_AX;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_A_CY;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_A_XOR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_B;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_B1;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_B2;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_B3;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_B4;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_B5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_B6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_BO5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_BO6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_B_CY;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_B_XOR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_C;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_C1;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_C2;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_C3;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_C4;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_C5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_C6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_CLK;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_CO5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_CO6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_C_CY;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_C_XOR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_D;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_D1;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_D2;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_D3;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_D4;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_D5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_D6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_DO5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_D_CY;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_D_XOR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X20Y152_SR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_A;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_A1;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_A2;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_A3;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_A4;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_A5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_A6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_AMUX;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_AO5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_AO6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_AQ;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_AX;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_A_CY;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_A_XOR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_B;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_B1;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_B2;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_B3;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_B4;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_B5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_B6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_BO5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_BO6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_BQ;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_BX;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_B_CY;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_B_XOR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_C;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_C1;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_C2;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_C3;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_C4;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_C5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_C6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_CLK;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_CMUX;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_CO5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_CO6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_C_CY;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_C_XOR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_D;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_D1;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_D2;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_D3;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_D4;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_D5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_D6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_DMUX;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_DO5;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_DO6;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_D_CY;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_D_XOR;
  wire [0:0] CLBLM_R_X15Y152_SLICE_X21Y152_SR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_AO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_AO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_BO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_BO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_CO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_CO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_DO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_DO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_AMUX;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_AO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_AO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_BO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_BO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_CMUX;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_CO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_CO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_DO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_DO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AMUX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CE;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CLK;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_SR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AQ;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BQ;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CLK;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_SR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CE;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_SR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_SR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CLK;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_SR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A5Q;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CLK;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_SR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CLK;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_DO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_DO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_SR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A5Q;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AMUX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CE;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CLK;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DMUX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_SR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CLK;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_SR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CE;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CLK;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_SR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CE;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CLK;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_SR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CLK;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_SR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CE;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CLK;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_SR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CLK;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_DMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_DO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_SR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CE;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CLK;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_COUT;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_SR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AMUX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CE;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CLK;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_SR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CE;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CIN;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CLK;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_COUT;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_SR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CLK;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_SR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CE;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CIN;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CLK;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_COUT;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_SR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CE;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CIN;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CLK;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_COUT;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_SR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CLK;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_SR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CLK;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_SR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CLK;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_SR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CLK;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_SR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CLK;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_SR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CLK;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_SR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AMUX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BMUX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CLK;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_SR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CE;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CLK;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_SR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CLK;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_SR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AQ;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CE;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CLK;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_SR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CLK;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_SR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AMUX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CE;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CLK;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_SR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CE;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CLK;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_SR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AQ;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AX;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_BO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CE;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CLK;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_DO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_SR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_BO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CLK;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_DO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_SR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A5Q;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AMUX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CE;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CLK;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CMUX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DMUX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_SR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CE;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CLK;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DQ;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_SR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AMUX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AQ;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_BO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_BQ;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_BX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CE;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CLK;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CQ;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_DO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_SR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_AQ;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_AX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_BO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_BO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_BQ;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_BX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CE;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CLK;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CQ;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_DO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_DO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_SR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CE;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CLK;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_SR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CE;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CLK;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DQ;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_SR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A5Q;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AMUX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CE;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CLK;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_SR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BMUX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CE;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CLK;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CMUX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DQ;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_SR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_A;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_A1;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_A2;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_A3;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_A4;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_A5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_A6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_AO5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_AO6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_AQ;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_AX;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_A_CY;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_A_XOR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_B;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_B1;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_B2;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_B3;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_B4;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_B5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_B6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_BO5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_BO6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_BQ;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_BX;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_B_CY;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_B_XOR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_C;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_C1;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_C2;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_C3;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_C4;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_C5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_C6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_CE;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_CLK;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_CO5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_CO6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_CQ;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_CX;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_C_CY;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_C_XOR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_D;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_D1;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_D2;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_D3;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_D4;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_D5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_D6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_DO5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_DO6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_DQ;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_DX;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_D_CY;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_D_XOR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X2Y159_SR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_A;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_A1;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_A2;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_A3;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_A4;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_A5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_A6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_AO5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_AO6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_AQ;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_AX;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_A_CY;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_A_XOR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_B;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_B1;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_B2;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_B3;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_B4;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_B5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_B6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_BO5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_BO6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_BQ;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_BX;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_B_CY;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_B_XOR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_C;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_C1;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_C2;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_C3;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_C4;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_C5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_C6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_CE;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_CLK;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_CO5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_CO6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_CQ;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_CX;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_C_CY;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_C_XOR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_D;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_D1;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_D2;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_D3;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_D4;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_D5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_D6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_DO5;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_DO6;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_D_CY;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_D_XOR;
  wire [0:0] CLBLM_R_X3Y159_SLICE_X3Y159_SR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CE;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_SR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_COUT;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CE;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_SR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CIN;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_COUT;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_COUT;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CIN;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_COUT;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CIN;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_COUT;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CIN;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_COUT;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CIN;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_COUT;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_SR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CIN;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_COUT;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CLK;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_SR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_SR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_SR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_SR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_SR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CLK;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_SR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CLK;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_SR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CLK;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_SR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CLK;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_SR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CLK;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_SR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CLK;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_SR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AMUX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CLK;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_SR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CE;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CLK;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_SR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CE;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CLK;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_SR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_F7AMUX_O;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_SR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CE;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_F7AMUX_O;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_SR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_COUT;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_F7AMUX_O;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CIN;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_COUT;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_F7AMUX_O;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CIN;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_COUT;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CLK;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_SR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_SR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CE;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_SR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CE;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CLK;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_SR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CE;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CLK;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_SR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CE;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_SR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CE;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_SR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CE;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_SR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_SR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_SR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CLK;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_SR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_SR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_F7AMUX_O;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_SR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_COUT;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CLK;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_SR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CIN;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_COUT;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_SR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CLK;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_F7AMUX_O;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_SR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_F7AMUX_O;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_SR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_SR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_SR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CE;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_SR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_SR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_SR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CLK;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_SR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_SR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CE;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_SR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_SR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CE;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_SR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CE;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_SR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CE;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CLK;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_SR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CE;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CLK;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_SR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CE;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_SR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_I;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_I;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_O;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_O;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_O;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_O;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_O;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_O;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_O;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_O;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_O;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_O;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_O;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_D;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_O;
  wire [0:0] LIOI3_SING_X0Y199_ILOGIC_X0Y199_D;
  wire [0:0] LIOI3_SING_X0Y199_ILOGIC_X0Y199_O;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_D1;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_OQ;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_T1;
  wire [0:0] LIOI3_SING_X0Y50_OLOGIC_X0Y50_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_O;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y167_D;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y167_O;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_D;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_O;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_D;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_O;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_D1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_OQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_T1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y51_TQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_D1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_OQ;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_T1;
  wire [0:0] LIOI3_X0Y51_OLOGIC_X0Y52_TQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_D1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_OQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_T1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y53_TQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_D1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_OQ;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_T1;
  wire [0:0] LIOI3_X0Y53_OLOGIC_X0Y54_TQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_D1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_OQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_T1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_TQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_D1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_OQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_T1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y56_TQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_D1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_OQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_T1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_TQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_D1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_OQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_T1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y60_TQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_D1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_OQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_T1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y61_TQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_D1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_OQ;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_T1;
  wire [0:0] LIOI3_X0Y61_OLOGIC_X0Y62_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_TQ;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_TQ;


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y116_SLICE_X0Y116_AO6),
.Q(CLBLL_L_X2Y116_SLICE_X0Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300330033003300)
  ) CLBLL_L_X2Y116_SLICE_X0Y116_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X0Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X0Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_DO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_CO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_BO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y116_SLICE_X1Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y116_SLICE_X1Y116_AO5),
.O6(CLBLL_L_X2Y116_SLICE_X1Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y132_SLICE_X2Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.Q(CLBLL_L_X2Y131_SLICE_X0Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y132_SLICE_X2Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_F7AMUX_O),
.Q(CLBLL_L_X2Y131_SLICE_X0Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I1(CLBLL_L_X2Y131_SLICE_X0Y131_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I5(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee000044440000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_BLUT (
.I0(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I1(CLBLL_L_X2Y131_SLICE_X0Y131_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc8c8cc44c840)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_ALUT (
.I0(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I2(CLBLL_L_X2Y131_SLICE_X0Y131_AQ),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I4(CLBLL_L_X2Y131_SLICE_X0Y131_BQ),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y132_SLICE_X2Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_DO6),
.Q(CLBLL_L_X2Y131_SLICE_X1Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_DO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_CO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_BO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_AO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y132_SLICE_X2Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.Q(CLBLL_L_X2Y132_SLICE_X1Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_DO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_CO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_BO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_AO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.Q(CLBLL_L_X2Y133_SLICE_X1Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_DO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_CO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_BO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X0Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X0Y135_AO5),
.O6(CLBLL_L_X2Y135_SLICE_X0Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y135_SLICE_X1Y135_AO5),
.Q(CLBLL_L_X2Y135_SLICE_X1Y135_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y135_SLICE_X1Y135_AO6),
.Q(CLBLL_L_X2Y135_SLICE_X1Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_DO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_CO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_BO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300330022222222)
  ) CLBLL_L_X2Y135_SLICE_X1Y135_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_CQ),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y135_SLICE_X1Y135_AO5),
.O6(CLBLL_L_X2Y135_SLICE_X1Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.Q(CLBLL_L_X2Y137_SLICE_X0Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.Q(CLBLL_L_X2Y137_SLICE_X0Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X0Y137_DO5),
.O6(CLBLL_L_X2Y137_SLICE_X0Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X0Y137_CO5),
.O6(CLBLL_L_X2Y137_SLICE_X0Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X0Y137_BO5),
.O6(CLBLL_L_X2Y137_SLICE_X0Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaccccff00)
  ) CLBLL_L_X2Y137_SLICE_X0Y137_ALUT (
.I0(CLBLL_L_X2Y138_SLICE_X0Y138_B_XOR),
.I1(CLBLL_L_X2Y137_SLICE_X0Y137_BQ),
.I2(CLBLL_L_X2Y137_SLICE_X0Y137_AQ),
.I3(CLBLL_L_X2Y138_SLICE_X0Y138_C_XOR),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X0Y137_AO5),
.O6(CLBLL_L_X2Y137_SLICE_X0Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X1Y137_DO5),
.O6(CLBLL_L_X2Y137_SLICE_X1Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X1Y137_CO5),
.O6(CLBLL_L_X2Y137_SLICE_X1Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afafa0a0)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_BLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_DQ),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I3(CLBLL_L_X2Y139_SLICE_X0Y139_B_XOR),
.I4(CLBLL_L_X2Y139_SLICE_X0Y139_C_XOR),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X1Y137_BO5),
.O6(CLBLL_L_X2Y137_SLICE_X1Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fafa0a0a)
  ) CLBLL_L_X2Y137_SLICE_X1Y137_ALUT (
.I0(CLBLL_L_X2Y139_SLICE_X0Y139_A_XOR),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I3(CLBLL_L_X2Y138_SLICE_X0Y138_D_XOR),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y137_SLICE_X1Y137_AO5),
.O6(CLBLL_L_X2Y137_SLICE_X1Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y138_SLICE_X0Y138_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X2Y138_SLICE_X0Y138_D_CY, CLBLL_L_X2Y138_SLICE_X0Y138_C_CY, CLBLL_L_X2Y138_SLICE_X0Y138_B_CY, CLBLL_L_X2Y138_SLICE_X0Y138_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLL_L_X2Y140_SLICE_X1Y140_BQ, 1'b0}),
.O({CLBLL_L_X2Y138_SLICE_X0Y138_D_XOR, CLBLL_L_X2Y138_SLICE_X0Y138_C_XOR, CLBLL_L_X2Y138_SLICE_X0Y138_B_XOR, CLBLL_L_X2Y138_SLICE_X0Y138_A_XOR}),
.S({CLBLL_L_X2Y138_SLICE_X0Y138_DO6, CLBLL_L_X2Y138_SLICE_X0Y138_CO6, CLBLL_L_X2Y138_SLICE_X0Y138_BO6, CLBLL_L_X2Y138_SLICE_X0Y138_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y140_SLICE_X1Y140_DQ),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y140_SLICE_X1Y140_CQ),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033007fffccff80)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I5(CLBLL_L_X2Y140_SLICE_X1Y140_BQ),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y140_SLICE_X1Y140_AQ),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y147_SLICE_X19Y147_BO6),
.Q(CLBLL_L_X2Y138_SLICE_X1Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y148_SLICE_X21Y148_BO6),
.Q(CLBLL_L_X2Y138_SLICE_X1Y138_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaccccff00)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_ALUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I1(CLBLL_L_X2Y138_SLICE_X1Y138_BQ),
.I2(CLBLL_L_X2Y138_SLICE_X1Y138_AQ),
.I3(CLBLL_L_X2Y138_SLICE_X0Y138_A_XOR),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y139_SLICE_X0Y139_CARRY4 (
.CI(CLBLL_L_X2Y138_SLICE_X0Y138_COUT),
.CO({CLBLL_L_X2Y139_SLICE_X0Y139_D_CY, CLBLL_L_X2Y139_SLICE_X0Y139_C_CY, CLBLL_L_X2Y139_SLICE_X0Y139_B_CY, CLBLL_L_X2Y139_SLICE_X0Y139_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X2Y139_SLICE_X0Y139_D_XOR, CLBLL_L_X2Y139_SLICE_X0Y139_C_XOR, CLBLL_L_X2Y139_SLICE_X0Y139_B_XOR, CLBLL_L_X2Y139_SLICE_X0Y139_A_XOR}),
.S({CLBLL_L_X2Y139_SLICE_X0Y139_DO6, CLBLL_L_X2Y139_SLICE_X0Y139_CO6, CLBLL_L_X2Y139_SLICE_X0Y139_BO6, CLBLL_L_X2Y139_SLICE_X0Y139_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y141_SLICE_X0Y141_AQ),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_DO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_CQ),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_CO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_BQ),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_BO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_AQ),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_AO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.Q(CLBLL_L_X2Y139_SLICE_X1Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.Q(CLBLL_L_X2Y139_SLICE_X1Y139_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.Q(CLBLL_L_X2Y139_SLICE_X1Y139_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_BO6),
.Q(CLBLL_L_X2Y139_SLICE_X1Y139_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50eeee4444)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I1(CLBLL_L_X2Y140_SLICE_X0Y140_A_XOR),
.I2(CLBLL_L_X2Y139_SLICE_X0Y139_D_XOR),
.I3(CLBLL_L_X2Y140_SLICE_X0Y140_BQ),
.I4(CLBLL_L_X2Y140_SLICE_X0Y140_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_DO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888f5a0f5a0)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_CLUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I1(CLBLL_L_X2Y139_SLICE_X1Y139_CQ),
.I2(CLBLL_L_X2Y139_SLICE_X1Y139_DQ),
.I3(CLBLL_L_X2Y141_SLICE_X0Y141_C_XOR),
.I4(CLBLL_L_X2Y141_SLICE_X0Y141_B_XOR),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_CO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccaaaa)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_BLUT (
.I0(CLBLL_L_X2Y141_SLICE_X0Y141_A_XOR),
.I1(CLBLL_L_X2Y139_SLICE_X1Y139_BQ),
.I2(CLBLL_L_X2Y140_SLICE_X0Y140_AQ),
.I3(CLBLL_L_X2Y140_SLICE_X0Y140_D_XOR),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_BO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_ALUT (
.I0(CLBLL_L_X2Y140_SLICE_X0Y140_B_XOR),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.I2(CLBLL_L_X2Y139_SLICE_X1Y139_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I4(CLBLL_L_X2Y140_SLICE_X0Y140_C_XOR),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_AO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y140_SLICE_X0Y140_AO5),
.Q(CLBLL_L_X2Y140_SLICE_X0Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y140_SLICE_X0Y140_BO5),
.Q(CLBLL_L_X2Y140_SLICE_X0Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y140_SLICE_X0Y140_CO5),
.Q(CLBLL_L_X2Y140_SLICE_X0Y140_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y140_SLICE_X0Y140_CARRY4 (
.CI(CLBLL_L_X2Y139_SLICE_X0Y139_COUT),
.CO({CLBLL_L_X2Y140_SLICE_X0Y140_D_CY, CLBLL_L_X2Y140_SLICE_X0Y140_C_CY, CLBLL_L_X2Y140_SLICE_X0Y140_B_CY, CLBLL_L_X2Y140_SLICE_X0Y140_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X2Y140_SLICE_X0Y140_D_XOR, CLBLL_L_X2Y140_SLICE_X0Y140_C_XOR, CLBLL_L_X2Y140_SLICE_X0Y140_B_XOR, CLBLL_L_X2Y140_SLICE_X0Y140_A_XOR}),
.S({CLBLL_L_X2Y140_SLICE_X0Y140_DO6, CLBLL_L_X2Y140_SLICE_X0Y140_CO6, CLBLL_L_X2Y140_SLICE_X0Y140_BO6, CLBLL_L_X2Y140_SLICE_X0Y140_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_DO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y143_SLICE_X1Y143_DQ),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_CO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00aaaaaaaa)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_BLUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X2Y142_SLICE_X1Y142_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_BO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_ALUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_BO6),
.I1(CLBLL_L_X2Y142_SLICE_X1Y142_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_AO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y140_SLICE_X1Y140_A_XOR),
.Q(CLBLL_L_X2Y140_SLICE_X1Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y140_SLICE_X1Y140_B_XOR),
.Q(CLBLL_L_X2Y140_SLICE_X1Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y140_SLICE_X1Y140_C_XOR),
.Q(CLBLL_L_X2Y140_SLICE_X1Y140_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y140_SLICE_X1Y140_D_XOR),
.Q(CLBLL_L_X2Y140_SLICE_X1Y140_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y140_SLICE_X1Y140_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X2Y140_SLICE_X1Y140_D_CY, CLBLL_L_X2Y140_SLICE_X1Y140_C_CY, CLBLL_L_X2Y140_SLICE_X1Y140_B_CY, CLBLL_L_X2Y140_SLICE_X1Y140_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLL_L_X2Y144_SLICE_X1Y144_CO6, 1'b0}),
.O({CLBLL_L_X2Y140_SLICE_X1Y140_D_XOR, CLBLL_L_X2Y140_SLICE_X1Y140_C_XOR, CLBLL_L_X2Y140_SLICE_X1Y140_B_XOR, CLBLL_L_X2Y140_SLICE_X1Y140_A_XOR}),
.S({CLBLL_L_X2Y140_SLICE_X1Y140_DO6, CLBLL_L_X2Y140_SLICE_X1Y140_CO6, CLBLL_L_X2Y140_SLICE_X1Y140_BO6, CLBLL_L_X2Y140_SLICE_X1Y140_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f1e0f5a0)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I2(CLBLL_L_X2Y140_SLICE_X1Y140_DQ),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_F7AMUX_O),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_DO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccccccaaa)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_CLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I1(CLBLL_L_X2Y140_SLICE_X1Y140_CQ),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_CO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666f66666660)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_BLUT (
.I0(CLBLL_L_X2Y144_SLICE_X1Y144_AO5),
.I1(CLBLL_L_X2Y140_SLICE_X1Y140_BQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_AO6),
.I5(CLBLL_L_X4Y141_SLICE_X4Y141_F7AMUX_O),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_BO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1f0e0f0f3f0c0)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I2(CLBLL_L_X2Y140_SLICE_X1Y140_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_F7AMUX_O),
.I5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_AO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y142_SLICE_X2Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y141_SLICE_X0Y141_AO5),
.Q(CLBLL_L_X2Y141_SLICE_X0Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y141_SLICE_X0Y141_CARRY4 (
.CI(CLBLL_L_X2Y140_SLICE_X0Y140_COUT),
.CO({CLBLL_L_X2Y141_SLICE_X0Y141_D_CY, CLBLL_L_X2Y141_SLICE_X0Y141_C_CY, CLBLL_L_X2Y141_SLICE_X0Y141_B_CY, CLBLL_L_X2Y141_SLICE_X0Y141_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X2Y141_SLICE_X0Y141_D_XOR, CLBLL_L_X2Y141_SLICE_X0Y141_C_XOR, CLBLL_L_X2Y141_SLICE_X0Y141_B_XOR, CLBLL_L_X2Y141_SLICE_X0Y141_A_XOR}),
.S({CLBLL_L_X2Y141_SLICE_X0Y141_DO6, CLBLL_L_X2Y141_SLICE_X0Y141_CO6, CLBLL_L_X2Y141_SLICE_X0Y141_BO6, CLBLL_L_X2Y141_SLICE_X0Y141_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_DO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y143_SLICE_X1Y143_CQ),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_CO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y143_SLICE_X1Y143_BQ),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_BO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y141_SLICE_X1Y141_D_XOR),
.I2(CLBLL_L_X2Y143_SLICE_X1Y143_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_AO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y141_SLICE_X1Y141_A_XOR),
.Q(CLBLL_L_X2Y141_SLICE_X1Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y141_SLICE_X1Y141_B_XOR),
.Q(CLBLL_L_X2Y141_SLICE_X1Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y141_SLICE_X1Y141_C_XOR),
.Q(CLBLL_L_X2Y141_SLICE_X1Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y141_SLICE_X1Y141_CARRY4 (
.CI(CLBLL_L_X2Y140_SLICE_X1Y140_COUT),
.CO({CLBLL_L_X2Y141_SLICE_X1Y141_D_CY, CLBLL_L_X2Y141_SLICE_X1Y141_C_CY, CLBLL_L_X2Y141_SLICE_X1Y141_B_CY, CLBLL_L_X2Y141_SLICE_X1Y141_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X2Y141_SLICE_X1Y141_D_XOR, CLBLL_L_X2Y141_SLICE_X1Y141_C_XOR, CLBLL_L_X2Y141_SLICE_X1Y141_B_XOR, CLBLL_L_X2Y141_SLICE_X1Y141_A_XOR}),
.S({CLBLL_L_X2Y141_SLICE_X1Y141_DO6, CLBLL_L_X2Y141_SLICE_X1Y141_CO6, CLBLL_L_X2Y141_SLICE_X1Y141_BO6, CLBLL_L_X2Y141_SLICE_X1Y141_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaba8bb88)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_DLUT (
.I0(CLBLL_L_X2Y141_SLICE_X0Y141_AQ),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_CO6),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_DO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fe04ee44)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_CLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_F7AMUX_O),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I3(CLBLL_L_X2Y141_SLICE_X1Y141_CQ),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_CO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccacccccaca)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_BLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_F7AMUX_O),
.I1(CLBLL_L_X2Y141_SLICE_X1Y141_BQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_BO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f0e4cc)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_F7AMUX_O),
.I2(CLBLL_L_X2Y141_SLICE_X1Y141_AQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_AO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y142_SLICE_X2Y142_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y142_SLICE_X1Y142_D_XOR),
.Q(CLBLL_L_X2Y142_SLICE_X0Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_DO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_CO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_BO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_AO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y142_SLICE_X2Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y142_SLICE_X1Y142_A_XOR),
.Q(CLBLL_L_X2Y142_SLICE_X1Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y142_SLICE_X2Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y142_SLICE_X1Y142_B_XOR),
.Q(CLBLL_L_X2Y142_SLICE_X1Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y142_SLICE_X1Y142_CARRY4 (
.CI(CLBLL_L_X2Y141_SLICE_X1Y141_COUT),
.CO({CLBLL_L_X2Y142_SLICE_X1Y142_D_CY, CLBLL_L_X2Y142_SLICE_X1Y142_C_CY, CLBLL_L_X2Y142_SLICE_X1Y142_B_CY, CLBLL_L_X2Y142_SLICE_X1Y142_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X2Y142_SLICE_X1Y142_D_XOR, CLBLL_L_X2Y142_SLICE_X1Y142_C_XOR, CLBLL_L_X2Y142_SLICE_X1Y142_B_XOR, CLBLL_L_X2Y142_SLICE_X1Y142_A_XOR}),
.S({CLBLL_L_X2Y142_SLICE_X1Y142_DO6, CLBLL_L_X2Y142_SLICE_X1Y142_CO6, CLBLL_L_X2Y142_SLICE_X1Y142_BO6, CLBLL_L_X2Y142_SLICE_X1Y142_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaabfaa80)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_DLUT (
.I0(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_CO6),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_DO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaba8afa0)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_CLUT (
.I0(CLBLL_L_X2Y143_SLICE_X1Y143_DQ),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_CO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccccdfcc80)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_BLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I1(CLBLL_L_X2Y142_SLICE_X1Y142_BQ),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_AO6),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_BO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1f0f3f0e0f0c0)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I2(CLBLL_L_X2Y142_SLICE_X1Y142_AQ),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I5(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_AO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y143_SLICE_X0Y143_AO6),
.Q(CLBLL_L_X2Y143_SLICE_X0Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_DO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_CO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_BO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0c0c0)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_AO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y142_SLICE_X2Y142_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y143_SLICE_X1Y143_A_XOR),
.Q(CLBLL_L_X2Y143_SLICE_X1Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y142_SLICE_X2Y142_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y143_SLICE_X1Y143_B_XOR),
.Q(CLBLL_L_X2Y143_SLICE_X1Y143_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y142_SLICE_X2Y142_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y143_SLICE_X1Y143_C_XOR),
.Q(CLBLL_L_X2Y143_SLICE_X1Y143_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y142_SLICE_X2Y142_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y143_SLICE_X1Y143_DO5),
.Q(CLBLL_L_X2Y143_SLICE_X1Y143_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y143_SLICE_X1Y143_CARRY4 (
.CI(CLBLL_L_X2Y142_SLICE_X1Y142_COUT),
.CO({CLBLL_L_X2Y143_SLICE_X1Y143_D_CY, CLBLL_L_X2Y143_SLICE_X1Y143_C_CY, CLBLL_L_X2Y143_SLICE_X1Y143_B_CY, CLBLL_L_X2Y143_SLICE_X1Y143_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X2Y143_SLICE_X1Y143_D_XOR, CLBLL_L_X2Y143_SLICE_X1Y143_C_XOR, CLBLL_L_X2Y143_SLICE_X1Y143_B_XOR, CLBLL_L_X2Y143_SLICE_X1Y143_A_XOR}),
.S({CLBLL_L_X2Y143_SLICE_X1Y143_DO6, CLBLL_L_X2Y143_SLICE_X1Y143_CO6, CLBLL_L_X2Y143_SLICE_X1Y143_BO6, CLBLL_L_X2Y143_SLICE_X1Y143_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_DLUT (
.I0(CLBLL_L_X2Y142_SLICE_X1Y142_C_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_DO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccccaccaa)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_CLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_AO6),
.I1(CLBLL_L_X2Y143_SLICE_X1Y143_CQ),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_CO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccdcfccccc8c0)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_BLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I1(CLBLL_L_X2Y143_SLICE_X1Y143_BQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_BO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0e4f0cc)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I1(CLBLM_R_X3Y144_SLICE_X3Y144_BO6),
.I2(CLBLL_L_X2Y143_SLICE_X1Y143_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_AO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y144_SLICE_X0Y144_AO5),
.Q(CLBLL_L_X2Y144_SLICE_X0Y144_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y144_SLICE_X0Y144_AO6),
.Q(CLBLL_L_X2Y144_SLICE_X0Y144_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_AO6),
.Q(CLBLL_L_X2Y144_SLICE_X0Y144_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_DO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_CO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_BO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_AO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_DO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff00ea00)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_CLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I3(CLBLL_L_X2Y144_SLICE_X1Y144_AO5),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_DO6),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_CO6),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_CO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c99fbff3933ffff)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_BLUT (
.I0(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_DO6),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I4(CLBLL_L_X2Y144_SLICE_X1Y144_AO6),
.I5(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_BO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f1f3fffffe0c0)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_ALUT (
.I0(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_AO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y145_SLICE_X0Y145_AO5),
.Q(CLBLL_L_X2Y145_SLICE_X0Y145_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y145_SLICE_X0Y145_AO6),
.Q(CLBLL_L_X2Y145_SLICE_X0Y145_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y145_SLICE_X1Y145_AO6),
.Q(CLBLL_L_X2Y145_SLICE_X1Y145_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffaaaaabaa)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I2(CLBLL_L_X2Y144_SLICE_X1Y144_BO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I5(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y147_SLICE_X0Y147_AO5),
.Q(CLBLL_L_X2Y147_SLICE_X0Y147_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.Q(CLBLL_L_X2Y147_SLICE_X0Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_ALUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLL_L_X2Y148_SLICE_X1Y148_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000a0a0a0a)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffefffe)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_BO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbcffbf01010101)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_DO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_CO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_BO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_AO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_DO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_CO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_BO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000011111100)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_ALUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_AO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y107_IOB_X0Y107_I),
.Q(CLBLL_L_X2Y152_SLICE_X0Y152_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_DO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_CO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_BO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_AO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_DO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_CO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_A5_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y107_IOB_X0Y107_I),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y193_IOB_X0Y194_I),
.Q(CLBLL_L_X2Y153_SLICE_X0Y153_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_B5_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y107_IOB_X0Y107_I),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y195_IOB_X0Y195_I),
.Q(CLBLL_L_X2Y153_SLICE_X0Y153_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_C5_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y107_IOB_X0Y107_I),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y195_IOB_X0Y196_I),
.Q(CLBLL_L_X2Y153_SLICE_X0Y153_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_D5_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y107_IOB_X0Y107_I),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y197_IOB_X0Y197_I),
.Q(CLBLL_L_X2Y153_SLICE_X0Y153_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y107_IOB_X0Y107_I),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y153_SLICE_X0Y153_AO6),
.Q(CLBLL_L_X2Y153_SLICE_X0Y153_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y107_IOB_X0Y107_I),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y153_SLICE_X0Y153_BO6),
.Q(CLBLL_L_X2Y153_SLICE_X0Y153_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y107_IOB_X0Y107_I),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y153_SLICE_X0Y153_CO6),
.Q(CLBLL_L_X2Y153_SLICE_X0Y153_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y107_IOB_X0Y107_I),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y153_SLICE_X0Y153_DO6),
.Q(CLBLL_L_X2Y153_SLICE_X0Y153_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y193_IOB_X0Y193_I),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_DO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y191_IOB_X0Y192_I),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_CO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y191_IOB_X0Y191_I),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_BO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y189_IOB_X0Y190_I),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_AO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y151_IOB_X0Y151_I),
.Q(CLBLL_L_X2Y153_SLICE_X1Y153_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y151_IOB_X0Y152_I),
.Q(CLBLL_L_X2Y153_SLICE_X1Y153_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00000000)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_DLUT (
.I0(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y153_SLICE_X0Y153_BQ),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_DO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ff55fa50aa00)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_CLUT (
.I0(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BQ),
.I3(CLBLL_L_X2Y153_SLICE_X0Y153_CQ),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I5(CLBLL_L_X2Y155_SLICE_X0Y155_BO6),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_CO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0f1f0f5f0f0f0)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_BLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_DO6),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_AO6),
.I5(CLBLM_R_X3Y156_SLICE_X3Y156_CO6),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_BO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0c0cff00d1d1)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_ALUT (
.I0(CLBLM_R_X3Y156_SLICE_X3Y156_CO6),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_AQ),
.I3(CLBLL_L_X2Y153_SLICE_X0Y153_BQ),
.I4(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y151_IOB_X0Y152_I),
.Q(CLBLL_L_X2Y155_SLICE_X0Y155_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y153_IOB_X0Y154_I),
.Q(CLBLL_L_X2Y155_SLICE_X0Y155_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_DO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfebafebafbfbeaea)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_CLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I2(CLBLL_L_X2Y158_SLICE_X1Y158_BQ),
.I3(CLBLL_L_X2Y155_SLICE_X0Y155_BQ),
.I4(CLBLL_L_X2Y157_SLICE_X0Y157_DO6),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_CO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3033300033220022)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_BLUT (
.I0(CLBLL_L_X2Y156_SLICE_X0Y156_DO6),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.I2(CLBLL_L_X2Y155_SLICE_X0Y155_AQ),
.I3(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I4(CLBLL_L_X2Y158_SLICE_X1Y158_AQ),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_BO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe1010ff00ff00)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_ALUT (
.I0(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I2(CLBLL_L_X2Y158_SLICE_X1Y158_AQ),
.I3(CLBLL_L_X2Y156_SLICE_X0Y156_AO6),
.I4(CLBLL_L_X2Y158_SLICE_X1Y158_DQ),
.I5(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_AO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y151_IOB_X0Y151_I),
.Q(CLBLL_L_X2Y155_SLICE_X1Y155_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_DO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_AO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y156_SLICE_X0Y156_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X1Y158_AQ),
.Q(CLBLL_L_X2Y156_SLICE_X0Y156_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y156_SLICE_X0Y156_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X1Y158_DQ),
.Q(CLBLL_L_X2Y156_SLICE_X0Y156_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y156_SLICE_X0Y156_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X0Y158_BQ),
.Q(CLBLL_L_X2Y156_SLICE_X0Y156_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y156_SLICE_X0Y156_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y155_SLICE_X0Y155_AQ),
.Q(CLBLL_L_X2Y156_SLICE_X0Y156_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffaaf0cc00aaf0)
  ) CLBLL_L_X2Y156_SLICE_X0Y156_DLUT (
.I0(CLBLL_L_X2Y156_SLICE_X0Y156_BQ),
.I1(CLBLL_L_X2Y156_SLICE_X0Y156_CQ),
.I2(CLBLL_L_X2Y156_SLICE_X0Y156_DQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLL_L_X2Y156_SLICE_X0Y156_AQ),
.O5(CLBLL_L_X2Y156_SLICE_X0Y156_DO5),
.O6(CLBLL_L_X2Y156_SLICE_X0Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafcfc0a0a0cfc0)
  ) CLBLL_L_X2Y156_SLICE_X0Y156_CLUT (
.I0(CLBLL_L_X2Y158_SLICE_X1Y158_AQ),
.I1(CLBLL_L_X2Y155_SLICE_X0Y155_AQ),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I3(CLBLL_L_X2Y156_SLICE_X0Y156_BQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLL_L_X2Y156_SLICE_X0Y156_CQ),
.O5(CLBLL_L_X2Y156_SLICE_X0Y156_CO5),
.O6(CLBLL_L_X2Y156_SLICE_X0Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fb73cc00c840)
  ) CLBLL_L_X2Y156_SLICE_X0Y156_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I2(CLBLL_L_X2Y158_SLICE_X1Y158_DQ),
.I3(CLBLL_L_X2Y158_SLICE_X0Y158_BQ),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I5(CLBLL_L_X2Y156_SLICE_X0Y156_CO6),
.O5(CLBLL_L_X2Y156_SLICE_X0Y156_BO5),
.O6(CLBLL_L_X2Y156_SLICE_X0Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdad5d0df8a85808)
  ) CLBLL_L_X2Y156_SLICE_X0Y156_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLL_L_X2Y156_SLICE_X0Y156_BQ),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I3(CLBLL_L_X2Y156_SLICE_X0Y156_CQ),
.I4(CLBLL_L_X2Y155_SLICE_X0Y155_AQ),
.I5(CLBLL_L_X2Y156_SLICE_X0Y156_AQ),
.O5(CLBLL_L_X2Y156_SLICE_X0Y156_AO5),
.O6(CLBLL_L_X2Y156_SLICE_X0Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y156_SLICE_X1Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y156_SLICE_X1Y156_DO5),
.O6(CLBLL_L_X2Y156_SLICE_X1Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y156_SLICE_X1Y156_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y156_SLICE_X1Y156_CO5),
.O6(CLBLL_L_X2Y156_SLICE_X1Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y156_SLICE_X1Y156_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y156_SLICE_X1Y156_BO5),
.O6(CLBLL_L_X2Y156_SLICE_X1Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y156_SLICE_X1Y156_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y156_SLICE_X1Y156_AO5),
.O6(CLBLL_L_X2Y156_SLICE_X1Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X1Y158_BQ),
.Q(CLBLL_L_X2Y157_SLICE_X0Y157_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X0Y158_AQ),
.Q(CLBLL_L_X2Y157_SLICE_X0Y157_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X0Y158_DQ),
.Q(CLBLL_L_X2Y157_SLICE_X0Y157_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y155_SLICE_X0Y155_BQ),
.Q(CLBLL_L_X2Y157_SLICE_X0Y157_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd8aad855d800d8)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLL_L_X2Y157_SLICE_X0Y157_AQ),
.I2(CLBLL_L_X2Y157_SLICE_X0Y157_DQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLL_L_X2Y157_SLICE_X0Y157_BQ),
.I5(CLBLL_L_X2Y157_SLICE_X0Y157_CQ),
.O5(CLBLL_L_X2Y157_SLICE_X0Y157_DO5),
.O6(CLBLL_L_X2Y157_SLICE_X0Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaddfa8850dd5088)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_CLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLL_L_X2Y157_SLICE_X0Y157_CQ),
.I2(CLBLL_L_X2Y155_SLICE_X0Y155_BQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLL_L_X2Y157_SLICE_X0Y157_BQ),
.I5(CLBLL_L_X2Y158_SLICE_X1Y158_BQ),
.O5(CLBLL_L_X2Y157_SLICE_X0Y157_CO5),
.O6(CLBLL_L_X2Y157_SLICE_X0Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_BLUT (
.I0(CLBLL_L_X2Y155_SLICE_X0Y155_BQ),
.I1(CLBLL_L_X2Y157_SLICE_X0Y157_BQ),
.I2(CLBLL_L_X2Y157_SLICE_X0Y157_AQ),
.I3(CLBLL_L_X2Y157_SLICE_X0Y157_CQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLL_L_X2Y157_SLICE_X0Y157_BO5),
.O6(CLBLL_L_X2Y157_SLICE_X0Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fc30aaaaaaaa)
  ) CLBLL_L_X2Y157_SLICE_X0Y157_ALUT (
.I0(CLBLL_L_X2Y157_SLICE_X0Y157_BO6),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I2(CLBLL_L_X2Y158_SLICE_X1Y158_BQ),
.I3(CLBLL_L_X2Y158_SLICE_X0Y158_AQ),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I5(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.O5(CLBLL_L_X2Y157_SLICE_X0Y157_AO5),
.O6(CLBLL_L_X2Y157_SLICE_X0Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X1Y157_DO5),
.O6(CLBLL_L_X2Y157_SLICE_X1Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X1Y157_CO5),
.O6(CLBLL_L_X2Y157_SLICE_X1Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X1Y157_BO5),
.O6(CLBLL_L_X2Y157_SLICE_X1Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y157_SLICE_X1Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y157_SLICE_X1Y157_AO5),
.O6(CLBLL_L_X2Y157_SLICE_X1Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_A5_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y179_IOB_X0Y180_I),
.Q(CLBLL_L_X2Y158_SLICE_X0Y158_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X0Y158_AO6),
.Q(CLBLL_L_X2Y158_SLICE_X0Y158_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y175_IOB_X0Y176_I),
.Q(CLBLL_L_X2Y158_SLICE_X0Y158_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y177_IOB_X0Y177_I),
.Q(CLBLL_L_X2Y158_SLICE_X0Y158_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y177_IOB_X0Y178_I),
.Q(CLBLL_L_X2Y158_SLICE_X0Y158_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X0Y158_DO5),
.O6(CLBLL_L_X2Y158_SLICE_X0Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X0Y158_CO5),
.O6(CLBLL_L_X2Y158_SLICE_X0Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fb73cc00c840)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_BLUT (
.I0(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I2(CLBLL_L_X2Y158_SLICE_X0Y158_AQ),
.I3(CLBLL_L_X2Y158_SLICE_X0Y158_DQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLL_L_X2Y157_SLICE_X0Y157_CO6),
.O5(CLBLL_L_X2Y158_SLICE_X0Y158_BO5),
.O6(CLBLL_L_X2Y158_SLICE_X0Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X2Y158_SLICE_X0Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y169_IOB_X0Y170_I),
.O5(CLBLL_L_X2Y158_SLICE_X0Y158_AO5),
.O6(CLBLL_L_X2Y158_SLICE_X0Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y159_IOB_X0Y160_I),
.Q(CLBLL_L_X2Y158_SLICE_X1Y158_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y161_IOB_X0Y162_I),
.Q(CLBLL_L_X2Y158_SLICE_X1Y158_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y163_IOB_X0Y164_I),
.Q(CLBLL_L_X2Y158_SLICE_X1Y158_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y167_IOB_X0Y168_I),
.Q(CLBLL_L_X2Y158_SLICE_X1Y158_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X1Y158_DO5),
.O6(CLBLL_L_X2Y158_SLICE_X1Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X1Y158_CO5),
.O6(CLBLL_L_X2Y158_SLICE_X1Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X1Y158_BO5),
.O6(CLBLL_L_X2Y158_SLICE_X1Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y158_SLICE_X1Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y158_SLICE_X1Y158_AO5),
.O6(CLBLL_L_X2Y158_SLICE_X1Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_AO5),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_AO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0dff08ff0dff08)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_DLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h40f0f000f000f000)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcddcddddcddccccc)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I5(CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0c3f0c2222eeee)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_ALUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_DO6),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_BO6),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fa00fafafafafa)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_ALUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y103_IOB_X0Y103_I),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111313111113131)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_ALUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_AO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_BO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2233222200330000)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I4(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fe00ccfefecccc)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I4(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5c5350ffcc3300)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_BLUT (
.I0(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5410febafc30fc30)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010ba101010ba10)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_DLUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_DO6),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_CO6),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h13335fff5fff5fff)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_CLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I5(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000eaaaffff)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_CO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.I5(CLBLL_L_X4Y134_SLICE_X5Y134_DO6),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cca0ec0000a0a0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddffff0ddd0fff)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_DLUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I5(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heac0c0c0aa000000)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_CLUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I5(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ffbfff)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I3(CLBLL_L_X4Y133_SLICE_X5Y133_DO6),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_DO6),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff5fff5fff0000)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_ALUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_AO6),
.I5(CLBLL_L_X4Y133_SLICE_X5Y133_CO6),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y133_SLICE_X5Y133_MUXF7A (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_AO6),
.O(CLBLL_L_X4Y133_SLICE_X5Y133_F7AMUX_O),
.S(CLBLM_R_X3Y133_SLICE_X3Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_BO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc00550005)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_DLUT (
.I0(LIOB33_SING_X0Y199_IOB_X0Y199_I),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.I4(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I5(CLBLM_R_X7Y135_SLICE_X8Y135_AO5),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ccc5fff4ccc4ccc)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_CLUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_DO6),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_AO5),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafaaaaafafaacc)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_DO6),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_AO5),
.I4(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.I5(CLBLM_R_X3Y134_SLICE_X2Y134_AO6),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c000000c0c0000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033113301)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_DO6),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_AO5),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_DO5),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ace00cc0a0a0000)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heccca000a000a000)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_BLUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c0c0c0c00000)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_AO5),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_BO5),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_CO5),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_DO5),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_AO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_BO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_CO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_DO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc0000ff00)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222fc30fc30)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.I3(CLBLM_R_X15Y139_SLICE_X21Y139_AO5),
.I4(CLBLM_R_X15Y141_SLICE_X20Y141_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505050ee44ee44)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_BLUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I1(CLBLM_R_X15Y140_SLICE_X21Y140_DO6),
.I2(CLBLM_R_X15Y142_SLICE_X20Y142_BO6),
.I3(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_AO5),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_BO5),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_CO5),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_AO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_BO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_CO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880000880088)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_DLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0aaf0aa)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.I2(CLBLM_R_X15Y140_SLICE_X21Y140_AO5),
.I3(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I4(CLBLM_R_X15Y143_SLICE_X21Y143_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h222222223300ffcc)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_DQ),
.I4(CLBLM_R_X13Y141_SLICE_X19Y141_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300330030303030)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y147_SLICE_X19Y147_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y148_SLICE_X21Y148_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000031000000)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h200030008000c000)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_BLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055aaff27272727)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(LIOB33_X0Y187_IOB_X0Y187_I),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I4(LIOB33_X0Y185_IOB_X0Y186_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd555d555c000c000)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_BLUT (
.I0(CLBLM_L_X10Y136_SLICE_X12Y136_CO6),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000300300030)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_AO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_CO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa50cccccccc)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.I2(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_BO5),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a2a2a2a2222aaaa)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_BLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf0d8f050f0d8)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_ALUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_AQ),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_BO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc8cdc8c8c8cdcdc)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f3333555500ff)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_ALUT (
.I0(LIOB33_X0Y185_IOB_X0Y185_I),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I2(LIOB33_X0Y183_IOB_X0Y183_I),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h080008000c000c00)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_BO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd800000072000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff50ff44cccccccc)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I1(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c04040c0ff40ff)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_ALUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_BO6),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I5(CLBLL_L_X4Y140_SLICE_X5Y140_CO6),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7c4f7f7f7c4c4c4)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_DLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_CO6),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I2(CLBLL_L_X4Y145_SLICE_X5Y145_AO6),
.I3(CLBLL_L_X4Y141_SLICE_X4Y141_CO6),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_BO6),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0aaaacccc)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR),
.I1(CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfb7373c8c84040)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_BLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR),
.I3(1'b1),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_AO6),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300ee22ee22)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y141_SLICE_X4Y141_MUXF7A (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_BO6),
.I1(CLBLL_L_X4Y141_SLICE_X4Y141_AO6),
.O(CLBLL_L_X4Y141_SLICE_X4Y141_F7AMUX_O),
.S(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y141_SLICE_X5Y141_AO5),
.Q(CLBLL_L_X4Y141_SLICE_X5Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.Q(CLBLL_L_X4Y141_SLICE_X5Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y141_SLICE_X5Y141_CO5),
.Q(CLBLL_L_X4Y141_SLICE_X5Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y141_SLICE_X5Y141_DO5),
.Q(CLBLL_L_X4Y141_SLICE_X5Y141_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X4Y141_SLICE_X5Y141_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X4Y141_SLICE_X5Y141_D_CY, CLBLL_L_X4Y141_SLICE_X5Y141_C_CY, CLBLL_L_X4Y141_SLICE_X5Y141_B_CY, CLBLL_L_X4Y141_SLICE_X5Y141_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X3Y140_SLICE_X3Y140_DQ, CLBLM_R_X3Y140_SLICE_X3Y140_CQ, CLBLM_R_X3Y140_SLICE_X3Y140_BQ, CLBLM_R_X3Y140_SLICE_X3Y140_AQ}),
.O({CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR, CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR, CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR, CLBLL_L_X4Y141_SLICE_X5Y141_A_XOR}),
.S({CLBLL_L_X4Y141_SLICE_X5Y141_DO6, CLBLL_L_X4Y141_SLICE_X5Y141_CO6, CLBLL_L_X4Y141_SLICE_X5Y141_BO6, CLBLL_L_X4Y141_SLICE_X5Y141_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf3003fcaaaaaaaa)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_BO6),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_BO6),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c333cccaaaaaaaa)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_CLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_BO6),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h772288ddf0f0f0f0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_BLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I3(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05affa50cccccccc)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_ALUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0f00000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR),
.I4(CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f4f7f7f0fcf3fff)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacaca00ff00ff)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_BLUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I3(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aafaccfacc)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_ALUT (
.I0(CLBLM_R_X15Y148_SLICE_X21Y148_BO6),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_DO6),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_L_X4Y142_SLICE_X4Y142_MUXF7A (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_AO6),
.O(CLBLL_L_X4Y142_SLICE_X4Y142_F7AMUX_O),
.S(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_BO5),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X4Y142_SLICE_X5Y142_CARRY4 (
.CI(CLBLL_L_X4Y141_SLICE_X5Y141_COUT),
.CO({CLBLL_L_X4Y142_SLICE_X5Y142_D_CY, CLBLL_L_X4Y142_SLICE_X5Y142_C_CY, CLBLL_L_X4Y142_SLICE_X5Y142_B_CY, CLBLL_L_X4Y142_SLICE_X5Y142_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X3Y141_SLICE_X3Y141_DQ, CLBLM_R_X3Y141_SLICE_X3Y141_CQ, CLBLM_R_X3Y141_SLICE_X3Y141_BQ, CLBLM_R_X3Y141_SLICE_X3Y141_AQ}),
.O({CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR, CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR, CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR, CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR}),
.S({CLBLL_L_X4Y142_SLICE_X5Y142_DO6, CLBLL_L_X4Y142_SLICE_X5Y142_CO6, CLBLL_L_X4Y142_SLICE_X5Y142_BO6, CLBLL_L_X4Y142_SLICE_X5Y142_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aaf0f0f0f0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_DO6),
.I3(CLBLM_R_X3Y141_SLICE_X3Y141_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa550ff0cccccccc)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_CO6),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_DO6),
.I3(CLBLM_R_X3Y141_SLICE_X3Y141_CQ),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66663c3cff00ff00)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.I1(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_CO6),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_AO6),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc0ff0aaaaaaaa)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_BO6),
.I3(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a500a500cc00cc)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_A_CY),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0c05f505f5)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.I1(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.I4(CLBLL_L_X4Y144_SLICE_X4Y144_CO6),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500500544444444)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_AO5),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_A_CY),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff50ff00ffcc)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.I2(CLBLM_R_X15Y148_SLICE_X21Y148_BO6),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_BO6),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X4Y143_SLICE_X5Y143_CARRY4 (
.CI(CLBLL_L_X4Y142_SLICE_X5Y142_COUT),
.CO({CLBLL_L_X4Y143_SLICE_X5Y143_D_CY, CLBLL_L_X4Y143_SLICE_X5Y143_C_CY, CLBLL_L_X4Y143_SLICE_X5Y143_B_CY, CLBLL_L_X4Y143_SLICE_X5Y143_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR, CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR, CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR, CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR}),
.S({CLBLL_L_X4Y143_SLICE_X5Y143_DO6, CLBLL_L_X4Y143_SLICE_X5Y143_CO6, CLBLL_L_X4Y143_SLICE_X5Y143_BO6, CLBLL_L_X4Y143_SLICE_X5Y143_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33ccf0f0f0f0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5aaa5aacccccccc)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0a5500ffaa5500)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_BLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I3(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I4(CLBLL_L_X2Y157_SLICE_X0Y157_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_ALUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_A_CY),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_AO5),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_BO5),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X4Y144_SLICE_X5Y144_CARRY4 (
.CI(CLBLL_L_X4Y143_SLICE_X5Y143_COUT),
.CO({CLBLL_L_X4Y144_SLICE_X5Y144_D_CY, CLBLL_L_X4Y144_SLICE_X5Y144_C_CY, CLBLL_L_X4Y144_SLICE_X5Y144_B_CY, CLBLL_L_X4Y144_SLICE_X5Y144_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR, CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR, CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR, CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR}),
.S({CLBLL_L_X4Y144_SLICE_X5Y144_DO6, CLBLL_L_X4Y144_SLICE_X5Y144_CO6, CLBLL_L_X4Y144_SLICE_X5Y144_BO6, CLBLL_L_X4Y144_SLICE_X5Y144_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000cccccccc)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4fcf4fcf40c040c0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_DLUT (
.I0(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_CO6),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5553333f5553333)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_CLUT (
.I0(CLBLL_L_X4Y155_SLICE_X4Y155_AO6),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccfcccccceeee)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.I1(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f552a00c0c0c0c0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_ALUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I3(CLBLL_L_X2Y156_SLICE_X0Y156_BO6),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h007700dd00220088)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_AO5),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_BO5),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0000e400)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I1(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I5(CLBLL_L_X4Y145_SLICE_X5Y145_BO6),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habaaabaaafaeabaa)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_DO6),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I2(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I4(CLBLM_R_X13Y147_SLICE_X19Y147_BO6),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00470047333333ff)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_ALUT (
.I0(CLBLM_L_X12Y146_SLICE_X16Y146_DO6),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00ccccff00cccc)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I3(CLBLL_L_X2Y155_SLICE_X0Y155_AO6),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff55550aaa0000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_BLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X3Y156_SLICE_X3Y156_AO6),
.I5(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbfbbffff)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_ALUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000c0000008c)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha08200880a080088)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_CLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_CO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff5f7f)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff75203030)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_BO6),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_AO6),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_AO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_DLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccccffffccee)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_CLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_DO6),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdcdcdcdcdcdd)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_BLUT (
.I0(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdcdcdcdddcdd)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_CO6),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_BO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100005555)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_DLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X5Y148_SLICE_X7Y148_BO5),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfffdccccccec)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_CLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_CO6),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_DO6),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_AO5),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_AO5),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddccddddddcc)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_BO6),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f03030a0a0000)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdfdedfffffffff)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_CO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff360000ffd60000)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050000018400000)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30300c0cf0f0feff)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_BO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080000800080)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_AO6),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000041000000)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f080f000f000f00)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_BLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BO6),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_AO5),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1155115533ff0000)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000d050f0f0f0f)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8105008091550080)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ee00ff00e000f0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_CO6),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.I4(CLBLL_L_X4Y149_SLICE_X4Y149_CO6),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_AO5),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa0000ffffeeee)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_DO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0c0cccec0cac)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_DLUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_BO5),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_BO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_BO6),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3fff3c3cc030c)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005533ef33ef)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4e020e02f7b316b2)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f0a0f050f0f)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_DLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00b100a000110000)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_CLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e0f000f0c0f000)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff80a2aaaa)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_BO6),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haffeaffffffefafa)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_DLUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd040500050505050)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffa000f2f2)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_CO6),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb00330033)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_DO5),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc33330f0f0f0f)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbfffffff3fff3)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_CLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I4(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000c0cffaaaeae)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_BLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_DO6),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_AO5),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_CO6),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14ff55ff55ee44)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_BO6),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000c000000100)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000200cc00ce00)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffaffbfffaffff)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbfbfaabbafbf)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_ALUT (
.I0(CLBLL_L_X4Y151_SLICE_X5Y151_DO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_DO6),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_BO6),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_CO5),
.I5(CLBLL_L_X4Y151_SLICE_X5Y151_CO6),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_DO5),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_DO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee222eeee22222)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_CLUT (
.I0(CLBLL_L_X4Y156_SLICE_X4Y156_BO6),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLL_L_X2Y158_SLICE_X0Y158_A5Q),
.I5(CLBLM_R_X3Y157_SLICE_X3Y157_BQ),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_CO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc88c8404400c840)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_BLUT (
.I0(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_BO6),
.I2(CLBLL_L_X4Y156_SLICE_X4Y156_AO6),
.I3(CLBLM_R_X3Y157_SLICE_X3Y157_BQ),
.I4(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I5(CLBLL_L_X2Y158_SLICE_X1Y158_CQ),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_BO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00efe04f40)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLM_R_X3Y159_SLICE_X3Y159_AQ),
.I2(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I3(CLBLM_R_X3Y155_SLICE_X3Y155_AO6),
.I4(CLBLM_R_X3Y159_SLICE_X2Y159_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_AO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_DO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_CO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_BO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_AO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X1Y158_CQ),
.Q(CLBLL_L_X4Y156_SLICE_X4Y156_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y157_SLICE_X3Y157_BQ),
.Q(CLBLL_L_X4Y156_SLICE_X4Y156_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X0Y158_A5Q),
.Q(CLBLL_L_X4Y156_SLICE_X4Y156_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y156_SLICE_X2Y156_AQ),
.Q(CLBLL_L_X4Y156_SLICE_X4Y156_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaccf000aaccf0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_DLUT (
.I0(CLBLL_L_X4Y156_SLICE_X4Y156_BQ),
.I1(CLBLL_L_X4Y156_SLICE_X4Y156_AQ),
.I2(CLBLL_L_X4Y156_SLICE_X4Y156_DQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I5(CLBLL_L_X4Y156_SLICE_X4Y156_CQ),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_DO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5550540405005404)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_CLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.I1(CLBLL_L_X4Y156_SLICE_X4Y156_DO6),
.I2(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.I3(CLBLL_L_X2Y158_SLICE_X1Y158_CQ),
.I4(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_AQ),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5ee44a0a0ee44)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLL_L_X4Y156_SLICE_X4Y156_BQ),
.I2(CLBLL_L_X2Y158_SLICE_X1Y158_CQ),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_CQ),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_AQ),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaad8d85500d8d8)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLL_L_X4Y156_SLICE_X4Y156_BQ),
.I2(CLBLL_L_X4Y156_SLICE_X4Y156_AQ),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_CQ),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_AQ),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_AO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_DO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_CO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_BO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_AO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303f3f05f505f5)
  ) CLBLL_L_X26Y133_SLICE_X38Y133_DLUT (
.I0(CLBLM_L_X16Y133_SLICE_X22Y133_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_L_X16Y133_SLICE_X23Y133_DQ),
.I5(1'b1),
.O5(CLBLL_L_X26Y133_SLICE_X38Y133_DO5),
.O6(CLBLL_L_X26Y133_SLICE_X38Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccaaaa)
  ) CLBLL_L_X26Y133_SLICE_X38Y133_CLUT (
.I0(CLBLM_L_X16Y134_SLICE_X23Y134_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X16Y133_SLICE_X23Y133_CQ),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I5(1'b1),
.O5(CLBLL_L_X26Y133_SLICE_X38Y133_CO5),
.O6(CLBLL_L_X26Y133_SLICE_X38Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055aaff1b1b1b1b)
  ) CLBLL_L_X26Y133_SLICE_X38Y133_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(CLBLM_L_X16Y133_SLICE_X22Y133_BQ),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X16Y133_SLICE_X23Y133_BQ),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLL_L_X26Y133_SLICE_X38Y133_BO5),
.O6(CLBLL_L_X26Y133_SLICE_X38Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44ee44)
  ) CLBLL_L_X26Y133_SLICE_X38Y133_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(CLBLM_L_X16Y133_SLICE_X22Y133_AQ),
.I2(CLBLM_L_X16Y133_SLICE_X23Y133_AQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X26Y133_SLICE_X38Y133_AO5),
.O6(CLBLL_L_X26Y133_SLICE_X38Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y133_SLICE_X39Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y133_SLICE_X39Y133_DO5),
.O6(CLBLL_L_X26Y133_SLICE_X39Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y133_SLICE_X39Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y133_SLICE_X39Y133_CO5),
.O6(CLBLL_L_X26Y133_SLICE_X39Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y133_SLICE_X39Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y133_SLICE_X39Y133_BO5),
.O6(CLBLL_L_X26Y133_SLICE_X39Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y133_SLICE_X39Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y133_SLICE_X39Y133_AO5),
.O6(CLBLL_L_X26Y133_SLICE_X39Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y135_SLICE_X38Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y135_SLICE_X38Y135_DO5),
.O6(CLBLL_L_X26Y135_SLICE_X38Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y135_SLICE_X38Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y135_SLICE_X38Y135_CO5),
.O6(CLBLL_L_X26Y135_SLICE_X38Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y135_SLICE_X38Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y135_SLICE_X38Y135_BO5),
.O6(CLBLL_L_X26Y135_SLICE_X38Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00e4e4e4e4)
  ) CLBLL_L_X26Y135_SLICE_X38Y135_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(CLBLM_L_X16Y135_SLICE_X22Y135_BQ),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_L_X16Y135_SLICE_X23Y135_AQ),
.I5(1'b1),
.O5(CLBLL_L_X26Y135_SLICE_X38Y135_AO5),
.O6(CLBLL_L_X26Y135_SLICE_X38Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y135_SLICE_X39Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y135_SLICE_X39Y135_DO5),
.O6(CLBLL_L_X26Y135_SLICE_X39Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y135_SLICE_X39Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y135_SLICE_X39Y135_CO5),
.O6(CLBLL_L_X26Y135_SLICE_X39Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y135_SLICE_X39Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y135_SLICE_X39Y135_BO5),
.O6(CLBLL_L_X26Y135_SLICE_X39Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y135_SLICE_X39Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y135_SLICE_X39Y135_AO5),
.O6(CLBLL_L_X26Y135_SLICE_X39Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X38Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X38Y136_DO5),
.O6(CLBLL_L_X26Y136_SLICE_X38Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X38Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X38Y136_CO5),
.O6(CLBLL_L_X26Y136_SLICE_X38Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00e4e4e4e4)
  ) CLBLL_L_X26Y136_SLICE_X38Y136_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(CLBLM_L_X16Y136_SLICE_X23Y136_CQ),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLM_L_X16Y136_SLICE_X23Y136_BQ),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X38Y136_BO5),
.O6(CLBLL_L_X26Y136_SLICE_X38Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505afaf22772277)
  ) CLBLL_L_X26Y136_SLICE_X38Y136_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(RIOB33_X105Y123_IOB_X1Y123_I),
.I2(CLBLM_L_X16Y136_SLICE_X23Y136_DQ),
.I3(CLBLM_L_X16Y139_SLICE_X22Y139_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X38Y136_AO5),
.O6(CLBLL_L_X26Y136_SLICE_X38Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X39Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X39Y136_DO5),
.O6(CLBLL_L_X26Y136_SLICE_X39Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X39Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X39Y136_CO5),
.O6(CLBLL_L_X26Y136_SLICE_X39Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X39Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X39Y136_BO5),
.O6(CLBLL_L_X26Y136_SLICE_X39Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X39Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X39Y136_AO5),
.O6(CLBLL_L_X26Y136_SLICE_X39Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y138_SLICE_X38Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y138_SLICE_X38Y138_DO5),
.O6(CLBLL_L_X26Y138_SLICE_X38Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y138_SLICE_X38Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y138_SLICE_X38Y138_CO5),
.O6(CLBLL_L_X26Y138_SLICE_X38Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y138_SLICE_X38Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y138_SLICE_X38Y138_BO5),
.O6(CLBLL_L_X26Y138_SLICE_X38Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLL_L_X26Y138_SLICE_X38Y138_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(RIOB33_X105Y115_IOB_X1Y115_I),
.I2(CLBLM_L_X16Y139_SLICE_X22Y139_AQ),
.I3(CLBLM_L_X16Y138_SLICE_X23Y138_AQ),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(1'b1),
.O5(CLBLL_L_X26Y138_SLICE_X38Y138_AO5),
.O6(CLBLL_L_X26Y138_SLICE_X38Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y138_SLICE_X39Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y138_SLICE_X39Y138_DO5),
.O6(CLBLL_L_X26Y138_SLICE_X39Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y138_SLICE_X39Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y138_SLICE_X39Y138_CO5),
.O6(CLBLL_L_X26Y138_SLICE_X39Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y138_SLICE_X39Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y138_SLICE_X39Y138_BO5),
.O6(CLBLL_L_X26Y138_SLICE_X39Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y138_SLICE_X39Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y138_SLICE_X39Y138_AO5),
.O6(CLBLL_L_X26Y138_SLICE_X39Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y101_IOB_X0Y102_I),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_BO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_CO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h050005000f0f0f0f)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_DO6),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055004400000044)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_CLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_DO6),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_AO6),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccccffffcccc)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccff0c0c0c0f)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff01ef0b4f)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_DLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0e0d0c0f1f2f3f)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010ffbf0013ffb3)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffb8b800fff0f0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I4(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b3ffffa0b3ffff)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_DLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I1(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.I2(LIOB33_SING_X0Y199_IOB_X0Y199_I),
.I3(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I4(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h437340704f7f4c7c)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_AO5),
.I4(CLBLL_L_X26Y133_SLICE_X38Y133_BO5),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5fffff00200000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_BLUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.I1(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333f0ff3333f000)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_BO6),
.I4(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef23e32cec20e02)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_DLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_BO6),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_BO6),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_AO6),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afafa0a0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_AO6),
.I1(CLBLM_L_X8Y135_SLICE_X11Y135_BO6),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_BO6),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_CO6),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fafa5050)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_BLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I1(CLBLM_R_X13Y136_SLICE_X19Y136_CO6),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_AO6),
.I3(CLBLM_L_X12Y134_SLICE_X16Y134_BO6),
.I4(CLBLM_R_X13Y133_SLICE_X19Y133_DO6),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44ee44)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_ALUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BO6),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_DO6),
.I4(CLBLM_L_X8Y133_SLICE_X10Y133_BO6),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X8Y134_SLICE_X10Y134_MUXF7A (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_BO6),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_AO6),
.O(CLBLM_L_X8Y134_SLICE_X10Y134_F7AMUX_O),
.S(CLBLM_R_X11Y143_SLICE_X14Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X8Y134_SLICE_X10Y134_MUXF7B (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_DO6),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_CO6),
.O(CLBLM_L_X8Y134_SLICE_X10Y134_F7BMUX_O),
.S(CLBLM_R_X11Y143_SLICE_X14Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X8Y134_SLICE_X10Y134_MUXF8 (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_F7BMUX_O),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_F7AMUX_O),
.O(CLBLM_L_X8Y134_SLICE_X10Y134_F8MUX_O),
.S(CLBLM_R_X7Y141_SLICE_X8Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050505050505050)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_DLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1b1b1b1b5500ffaa)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_CLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_CO5),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.I3(CLBLL_L_X26Y133_SLICE_X38Y133_BO6),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h01fb00ff01fb03f3)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ee00fc11ff03ff)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_ALUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I3(CLBLM_L_X16Y136_SLICE_X22Y136_BQ),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_AQ),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_BO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h505f505f30303f3f)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_DLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff05f511dd)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_CLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I1(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0e04fcfcfef4)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.I5(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f0dd11)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_ALUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000000000000)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000200000000000)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00030101ffcfefef)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_BLUT (
.I0(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2c0e2f3f0c0f0f3)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.I2(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I5(CLBLM_L_X8Y135_SLICE_X11Y135_CO6),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y136_SLICE_X10Y136_AO6),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y136_SLICE_X10Y136_BO6),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e2e2f0e2f0e2)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_AO5),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_AO6),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505050f7ffffff)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I2(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_BO6),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c5f5c505c5c5c5c)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_BLUT (
.I0(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_AO5),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0fad850d8)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_ALUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I5(CLBLM_L_X12Y137_SLICE_X16Y137_CO6),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y136_SLICE_X11Y136_AO6),
.Q(CLBLM_L_X8Y136_SLICE_X11Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f3f3f3f3)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000004000)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_DO6),
.I5(CLBLM_L_X8Y136_SLICE_X11Y136_BO6),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaf00550000)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4b0f4b0b0b0f4)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_ALUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_BO6),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_BO6),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaf0aa0faaff)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_CO6),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_AO5),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f5f305f3f503050)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_AO5),
.I1(CLBLM_L_X16Y137_SLICE_X23Y137_AO5),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I5(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacfcccccac0cccc)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_AO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I5(CLBLM_R_X15Y148_SLICE_X21Y148_BO6),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_DO6),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.I4(CLBLM_L_X8Y137_SLICE_X10Y137_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_AO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_BO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88ddfafa88dd5050)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(CLBLM_L_X16Y137_SLICE_X22Y137_AO5),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000000088000000)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_CLUT (
.I0(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdc8c8cdc8c8c)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_BLUT (
.I0(CLBLM_L_X12Y137_SLICE_X16Y137_CO5),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heef0f0f022f0f0f0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_ALUT (
.I0(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_BO6),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffaaaaaaaa)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_DLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7474747400ff00ff)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_CLUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(CLBLL_L_X26Y136_SLICE_X38Y136_AO6),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc747433ff)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.I3(CLBLM_R_X15Y140_SLICE_X21Y140_AO5),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000004e4e5f0a)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_R_X15Y142_SLICE_X20Y142_BO6),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f55550a0a0000)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_DLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7f7f5fff5f5f)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2fff2fffffff2fff)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_AO5),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff73ff7fc000c000)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_DO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333b7777777f)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_BO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_CO6),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_BO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c080c000000000)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_CLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_DO6),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_DO6),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff0fff11ff0fff)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_BO6),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_BO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_CO6),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000030377007700)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_ALUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_AO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4ccf5ffc4ccf5ff)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaeaaaaaaaaaaaa)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_AO6),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I5(CLBLM_L_X10Y136_SLICE_X12Y136_BO6),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffffff)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_DO6),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AO6),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I4(CLBLM_L_X8Y141_SLICE_X11Y141_AO6),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf80ff000a0a0000)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_BO6),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I3(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h005500550f0f0f0f)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_BO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff3300550055)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0e00000f000)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AO6),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_AO6),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbfff0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_ALUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_AO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c03c0300c03c030)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_BO6),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_AO5),
.I4(CLBLM_L_X8Y138_SLICE_X11Y138_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AO6),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f00008800)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I4(CLBLM_L_X8Y140_SLICE_X11Y140_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff00eeeef0f0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_ALUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_DO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f4f0f00004400)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_DLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_BO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLL_L_X4Y141_SLICE_X5Y141_DQ),
.I5(CLBLM_R_X5Y140_SLICE_X6Y140_BO6),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33113f153f153f15)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I2(CLBLM_R_X5Y148_SLICE_X7Y148_CO6),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2323afafff003333)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_DO6),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f500f5f5)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_ALUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_DO6),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0800070f00000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I3(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.I4(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4eeee4444444)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_AO5),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a00000fd08ff00)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_BO6),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_BO6),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d2e1d2ed1e2d1e2)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_DLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_AO6),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef2fe020afafa0a0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I1(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf870f870ffff0000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffa2aad5558000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y141_SLICE_X20Y141_DO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_AO5),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fffc0f000f0c)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_CO6),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_BO6),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha55a5aa55aa5a55a)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_AO5),
.I1(1'b1),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_AO5),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee22eaeeee222a)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_BLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_A5Q),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff20ff20df00df00)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3caaaa0f0f5555)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AO6),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_BO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h04c437f744447777)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaafbbbbfaffbbbb)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I1(CLBLM_R_X13Y147_SLICE_X19Y147_BO6),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AO6),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2aaaaff00ff00)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_R_X15Y148_SLICE_X21Y148_BO6),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafc0c0a0afc0c)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_DLUT (
.I0(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_BO6),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_DQ),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffacf0ac0fac00ac)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_CLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_CO6),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080000000800000)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc99c63366336c99c)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_ALUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_BO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_BO6),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0c0c0c0c)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heef5eea044f544a0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5353535300f00fff)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_CLUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00330f55ff330f55)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_DO6),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I2(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc4c4c4c40c040800)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fffffff5ffffff)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_CQ),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_DO6),
.I3(CLBLM_L_X8Y145_SLICE_X10Y145_AO5),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_AO6),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0fffffff7777)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_CLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_CQ),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_DO6),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50665033af66af33)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_BLUT (
.I0(CLBLM_R_X11Y145_SLICE_X14Y145_DO6),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_CQ),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_ALUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h001b551baa1bff1b)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_DLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I4(CLBLM_R_X3Y141_SLICE_X3Y141_DQ),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f75073fdffdcff)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_CLUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f0f7f0f0f0fff0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_BO6),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_AO6),
.I3(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30fcfc3074b874b8)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_ALUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_AO6),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f005f555faa5fff)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h11aa11ffbbaabbff)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_BO6),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0fff0dfc0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I4(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaefffbaff)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_BLUT (
.I0(CLBLM_R_X11Y147_SLICE_X15Y147_CO6),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_DO6),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_AO5),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I4(CLBLM_R_X7Y145_SLICE_X9Y145_DO6),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_CO6),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h007700f500dd00f5)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_ALUT (
.I0(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_DO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_BO6),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_AO5),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff7feeee)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd3c6c7c7d7d6d7d7)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00080f0f00080f0f)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_BO6),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f11bb5f5f11bb)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_BLUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_CO6),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000082000000ffff)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X15Y143_SLICE_X20Y143_AO5),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_F7AMUX_O),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555522222222)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_ALUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_BO6),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000039330000b9b3)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdecfd442200aa)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_CLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000200000002ff)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_L_X16Y142_SLICE_X22Y142_AO5),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_BO5),
.I3(CLBLM_L_X8Y149_SLICE_X10Y149_DO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I5(CLBLM_L_X8Y149_SLICE_X10Y149_CO6),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff9c0400000088)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_ALUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hec606cacff7f7fbf)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcff3cfffcfffcfff)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_AO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X8Y149_SLICE_X11Y149_MUXF7A (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_BO6),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_AO6),
.O(CLBLM_L_X8Y149_SLICE_X11Y149_F7AMUX_O),
.S(CLBLM_R_X3Y152_SLICE_X2Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101000011334444)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aa004d008800)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfffbfff3ffd3ff)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_BLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcececfcfcecececf)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_DO6),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_CO5),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_CO6),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000f58a8a00a0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcafacacafafafafa)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_BLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_AO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff05ff07ff05ff05)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_BO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_CO5),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb7bbbbb7b7bbbbb)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_BLUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I1(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I5(CLBLM_L_X12Y130_SLICE_X17Y130_BO6),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9333333380000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I1(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080008000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_CLUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I1(CLBLM_L_X12Y130_SLICE_X17Y130_BO6),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ceec0ee0)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I1(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.I5(CLBLM_L_X10Y130_SLICE_X13Y130_CO6),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h880000008f0f0f0f)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_ALUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I1(CLBLM_L_X12Y130_SLICE_X17Y130_BO6),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff30303030)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33b33333fff5ffff)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.I2(CLBLM_L_X12Y132_SLICE_X17Y132_B5Q),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff02ff0aff)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I5(CLBLM_L_X10Y131_SLICE_X12Y131_CO6),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haf8fa080af0fa000)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_BO6),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5ff80aaffd5aa80)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_DLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffba55005510)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_DO6),
.I4(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb8b8b8b8b8b8b8b)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_ALUT (
.I0(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I3(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fdddeccc)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_DO6),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00a0ffb3ff)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3fffff0faf0f8)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_DO6),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.I4(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00d800f0005000f0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_BO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_A5Q),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0c0c0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_B5Q),
.I2(CLBLM_L_X12Y132_SLICE_X17Y132_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h51fbfb5140eaea40)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_A5Q),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I5(CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00caca00000f0f)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_A_CY),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_D_CY),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I4(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500ffaacccccccc)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_CLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y131_SLICE_X18Y131_AO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff00f0cccccccc)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I3(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_AO6),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f0aaf033f0aaf0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I1(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacaff0ff000)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_ALUT (
.I0(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h500350f35f035ff3)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_CLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I1(CLBLL_L_X26Y133_SLICE_X38Y133_AO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e1f0c3f0e1f)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_BLUT (
.I0(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aa33f0f0f0f0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_DO6),
.I5(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h550f550f33ff3300)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I4(CLBLL_L_X26Y133_SLICE_X38Y133_DO6),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5c0c00000)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_BO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_CO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0530f530053ff53f)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_DLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf5a0dd88)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_CLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_DO6),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccaccc0cccacccf)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_AO6),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcfffdffff)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000200)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h437340704f7f4c7c)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_CLUT (
.I0(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.I4(CLBLL_L_X26Y133_SLICE_X38Y133_DO5),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000020003fffffff)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_BLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111000000003000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_AO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc00cc00cc)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffaaaaffff)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_CLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc0000fffff0f0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5b1b1e4e4a0a0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_DO6),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AO6),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff2fffffff)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_DLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_CLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_BO5),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_DO6),
.I5(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfdfd0c0c0000)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_BLUT (
.I0(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.I3(1'b1),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f0f0f00a0a0a0a)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_ALUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I1(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_BO6),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_CO6),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fe02aea2)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_AO6),
.I1(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccd8ccd8cc88ccdd)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_CLUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_L_X12Y137_SLICE_X16Y137_CO5),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccccccaa0f)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I2(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.I5(CLBLM_L_X12Y137_SLICE_X16Y137_CO6),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33553355000fff0f)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_ALUT (
.I0(CLBLM_R_X13Y138_SLICE_X19Y138_AQ),
.I1(RIOB33_X105Y115_IOB_X1Y116_I),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I4(LIOB33_X0Y187_IOB_X0Y188_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y137_SLICE_X13Y137_AO6),
.Q(CLBLM_L_X10Y137_SLICE_X13Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y137_SLICE_X13Y137_BO6),
.Q(CLBLM_L_X10Y137_SLICE_X13Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y137_SLICE_X13Y137_CO6),
.Q(CLBLM_L_X10Y137_SLICE_X13Y137_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y137_SLICE_X13Y137_DO6),
.Q(CLBLM_L_X10Y137_SLICE_X13Y137_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa3aca0afa3aca0)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_DLUT (
.I0(CLBLM_R_X13Y147_SLICE_X19Y147_BO6),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.I3(CLBLM_R_X13Y135_SLICE_X18Y135_BO6),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0efe0ef202f202)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_CLUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_AO6),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_DO6),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54ae04ae04)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_DO6),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I3(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.I4(1'b1),
.I5(CLBLM_R_X13Y137_SLICE_X18Y137_DO6),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fa50af05aa00)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.I1(1'b1),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I3(CLBLM_R_X15Y148_SLICE_X21Y148_BO6),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_AO6),
.I5(CLBLM_L_X12Y135_SLICE_X17Y135_DO6),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0fff08888bbbb)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_DLUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I2(CLBLM_R_X15Y138_SLICE_X21Y138_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff5500c5c5c5c5)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_CLUT (
.I0(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.I4(CLBLM_R_X15Y137_SLICE_X21Y137_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8008000055000000)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_AO6),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaad0d0dddd)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_DO6),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_AO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y138_SLICE_X13Y138_AO6),
.Q(CLBLM_L_X10Y138_SLICE_X13Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_BLUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_AO6),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_AO5),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacacfc0cfc0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_ALUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_CO6),
.I1(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_AO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.Q(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X12Y139_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X10Y139_SLICE_X12Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.Q(CLBLM_L_X10Y139_SLICE_X12Y139_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000033330000a55a)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_AO6),
.I1(CLBLM_R_X13Y131_SLICE_X18Y131_AQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaf0f0f033f0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X15Y144_SLICE_X21Y144_CO6),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_DO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb000b0fff000f0ff)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_CLUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_CO6),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00008000)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I5(CLBLM_L_X10Y139_SLICE_X13Y139_CO6),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccceefecccceeff)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_ALUT (
.I0(CLBLM_L_X12Y139_SLICE_X17Y139_CO6),
.I1(CLBLM_R_X11Y137_SLICE_X15Y137_AO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X11Y135_SLICE_X15Y135_AO5),
.I4(CLBLM_R_X11Y138_SLICE_X15Y138_BO6),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_CO6),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2233223322332233)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_CLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdfcfffccffccff)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a008a002000aa00)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_AO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_BO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044337700443377)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000088084404)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_CLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_AO5),
.I2(CLBLM_L_X12Y138_SLICE_X17Y138_BO6),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_CO6),
.I4(CLBLM_L_X8Y140_SLICE_X11Y140_AO6),
.I5(CLBLM_R_X13Y140_SLICE_X19Y140_BO6),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd5df858ad0da808)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_BO6),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.I4(CLBLM_L_X12Y142_SLICE_X16Y142_BO6),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cfcfc0c0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_ALUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_AO6),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_AO6),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.I3(CLBLM_R_X11Y141_SLICE_X14Y141_AO6),
.I4(CLBLM_L_X12Y142_SLICE_X16Y142_AO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_AO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AO5),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff7777ff)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_CLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_CO6),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AO5),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_DO6),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_BO6),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9ff9ffff9ff99ff9)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_BO5),
.I1(CLBLM_R_X11Y138_SLICE_X15Y138_DO6),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_DO6),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_CO6),
.I4(CLBLM_L_X12Y138_SLICE_X17Y138_BO6),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_CO6),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000000c00000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_DO6),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_DO6),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_BO6),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_CO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AO5),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfa0afa0a)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_DLUT (
.I0(CLBLM_R_X15Y148_SLICE_X21Y148_BO6),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_DO6),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff0013005f)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AO6),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I5(CLBLM_R_X11Y146_SLICE_X15Y146_AO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc693396c396cc693)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00f3f333f3)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y142_SLICE_X17Y142_DO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_BO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fedcfa503210)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_DLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I4(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I5(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0efec2320)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I5(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeef0fcaa22f030)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_BLUT (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.I3(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(CLBLM_L_X10Y137_SLICE_X13Y137_DQ),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff55550f0f)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_BO6),
.I3(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fafa5050)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_CLUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefc302222fc30)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_BLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_CO6),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_CQ),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h11110a5fbbbb0a5f)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc0000cccc)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11ddcfcf11ddcfcf)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_DO6),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd5da808fc0cfc0c)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_BLUT (
.I0(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_CQ),
.I4(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.I5(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h003305ff0033afff)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.I2(CLBLM_R_X11Y142_SLICE_X15Y142_F8MUX_O),
.I3(CLBLM_L_X8Y149_SLICE_X10Y149_BQ),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X10Y144_SLICE_X12Y144_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X10Y144_SLICE_X12Y144_D_CY, CLBLM_L_X10Y144_SLICE_X12Y144_C_CY, CLBLM_L_X10Y144_SLICE_X12Y144_B_CY, CLBLM_L_X10Y144_SLICE_X12Y144_A_CY}),
.CYINIT(CLBLM_L_X12Y144_SLICE_X16Y144_DO6),
.DI({CLBLM_R_X11Y144_SLICE_X15Y144_AO6, CLBLM_R_X11Y144_SLICE_X14Y144_DO6, CLBLM_L_X10Y144_SLICE_X13Y144_DO6, CLBLM_L_X10Y144_SLICE_X12Y144_AO5}),
.O({CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR, CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR, CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR, CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR}),
.S({CLBLM_L_X10Y144_SLICE_X12Y144_DO6, CLBLM_L_X10Y144_SLICE_X12Y144_CO6, CLBLM_L_X10Y144_SLICE_X12Y144_BO6, CLBLM_L_X10Y144_SLICE_X12Y144_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05af05af22227777)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_DLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I2(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_DO6),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2700275527aa27ff)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff333355550f0f)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_BLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0033333333)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333300ff00ff)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0bab0bab5bfb5bfb)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_CO6),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffddffcf)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_BLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccefccec)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X10Y145_SLICE_X12Y145_CARRY4 (
.CI(CLBLM_L_X10Y144_SLICE_X12Y144_COUT),
.CO({CLBLM_L_X10Y145_SLICE_X12Y145_D_CY, CLBLM_L_X10Y145_SLICE_X12Y145_C_CY, CLBLM_L_X10Y145_SLICE_X12Y145_B_CY, CLBLM_L_X10Y145_SLICE_X12Y145_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X10Y145_SLICE_X13Y145_DO6, CLBLM_R_X11Y145_SLICE_X15Y145_CO6, CLBLM_L_X10Y144_SLICE_X13Y144_DO5, CLBLM_L_X10Y145_SLICE_X13Y145_DO5}),
.O({CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR, CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR, CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR, CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR}),
.S({CLBLM_L_X10Y145_SLICE_X12Y145_DO6, CLBLM_L_X10Y145_SLICE_X12Y145_CO6, CLBLM_L_X10Y145_SLICE_X12Y145_BO6, CLBLM_L_X10Y145_SLICE_X12Y145_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505afafbbbbbbbb)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I5(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h220a770a225f775f)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I4(CLBLM_R_X3Y141_SLICE_X3Y141_DQ),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555505115555)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_BLUT (
.I0(CLBLM_R_X7Y145_SLICE_X9Y145_BO6),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I2(CLBLM_R_X3Y141_SLICE_X3Y141_CQ),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h404c707c434f737f)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I3(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_CO6),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff55555555)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a3b6e7f2a3b6e7f)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000afbfffbf)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_BLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I4(CLBLM_R_X3Y141_SLICE_X3Y141_CQ),
.I5(CLBLM_R_X7Y145_SLICE_X9Y145_BO6),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h550f3300550f33ff)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I1(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_CO6),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X10Y146_SLICE_X12Y146_CARRY4 (
.CI(CLBLM_L_X10Y145_SLICE_X12Y145_COUT),
.CO({CLBLM_L_X10Y146_SLICE_X12Y146_D_CY, CLBLM_L_X10Y146_SLICE_X12Y146_C_CY, CLBLM_L_X10Y146_SLICE_X12Y146_B_CY, CLBLM_L_X10Y146_SLICE_X12Y146_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X10Y147_SLICE_X13Y147_DO6, CLBLM_L_X10Y147_SLICE_X13Y147_DO5, CLBLM_L_X10Y148_SLICE_X12Y148_DO6, CLBLM_R_X11Y147_SLICE_X14Y147_DO6}),
.O({CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR, CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR, CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR, CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR}),
.S({CLBLM_L_X10Y146_SLICE_X12Y146_DO6, CLBLM_L_X10Y146_SLICE_X12Y146_CO6, CLBLM_L_X10Y146_SLICE_X12Y146_BO6, CLBLM_L_X10Y146_SLICE_X12Y146_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505bbbbafafbbbb)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_BO6),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2727aaff2727aaff)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_CO6),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff000f55ffff0f)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff0a0a55ff5f5f)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_DO6),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0bab0bab5bfb5bfb)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf00cf008b00cf00)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I2(CLBLM_L_X12Y143_SLICE_X16Y143_BO5),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc3ff55ff00ff00)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_CO6),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_AO6),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd11dd1d100000000)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_AO6),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_BO6),
.I4(CLBLM_L_X8Y145_SLICE_X10Y145_AO5),
.I5(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X10Y147_SLICE_X12Y147_CARRY4 (
.CI(CLBLM_L_X10Y146_SLICE_X12Y146_COUT),
.CO({CLBLM_L_X10Y147_SLICE_X12Y147_D_CY, CLBLM_L_X10Y147_SLICE_X12Y147_C_CY, CLBLM_L_X10Y147_SLICE_X12Y147_B_CY, CLBLM_L_X10Y147_SLICE_X12Y147_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLM_L_X10Y148_SLICE_X13Y148_DO6, CLBLM_R_X11Y147_SLICE_X14Y147_DO5}),
.O({CLBLM_L_X10Y147_SLICE_X12Y147_D_XOR, CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR, CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR, CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR}),
.S({CLBLM_L_X10Y147_SLICE_X12Y147_DO6, CLBLM_L_X10Y147_SLICE_X12Y147_CO6, CLBLM_L_X10Y147_SLICE_X12Y147_BO6, CLBLM_L_X10Y147_SLICE_X12Y147_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a2a2f2f7a7a7f7f)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y143_SLICE_X15Y143_CO6),
.I5(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55551b1bffff1b1b)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_BLUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_BO6),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I5(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff0f33ffff0f33)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f33333333)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff53a3ffff0000)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_CLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_BO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_AO5),
.I4(CLBLM_L_X12Y146_SLICE_X17Y146_F7AMUX_O),
.I5(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffff)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AO6),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_BO6),
.I2(CLBLM_L_X8Y145_SLICE_X10Y145_AO6),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.I4(CLBLM_R_X7Y145_SLICE_X9Y145_AO6),
.I5(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfff4fff2222bbbb)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_ALUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_BO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a200a2aaa20aa2)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_CLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_AO6),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_BO6),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_DO6),
.I5(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdf7757ffffffff)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333aaaa0f0f)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_ALUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I1(CLBLM_R_X13Y147_SLICE_X18Y147_C_XOR),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e200cc33ff)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I3(CLBLM_R_X13Y147_SLICE_X18Y147_B_XOR),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7f3f3fff7f)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_CO6),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00e000e0eaeaeaea)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_BQ),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I3(CLBLM_R_X11Y143_SLICE_X15Y143_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeffffdeeffdfdef)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_BO6),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7effe7ff9ffff9)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffb7edffffdb7e)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_CLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_DO6),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffdffdf7df)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_AO5),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I5(CLBLM_L_X10Y149_SLICE_X13Y149_CO6),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0517ffff175fffff)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_BO6),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h010007051f0f7f5f)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(CLBLM_R_X15Y150_SLICE_X21Y150_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AO6),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8cef08ce5a5a5a5a)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I4(CLBLM_R_X11Y150_SLICE_X15Y150_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff17055f17)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_BO6),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(CLBLM_R_X15Y151_SLICE_X20Y151_BO6),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a17055f17)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_BO6),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y128_SLICE_X16Y128_BO6),
.D(CLBLM_L_X12Y128_SLICE_X16Y128_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X12Y128_SLICE_X16Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050504000505)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_AO6),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_BO6),
.I4(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I5(CLBLM_R_X13Y128_SLICE_X18Y128_CO6),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddfffffcffffff)
  ) CLBLM_L_X12Y128_SLICE_X16Y128_ALUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I1(CLBLM_R_X15Y129_SLICE_X21Y129_BQ),
.I2(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I4(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I5(CLBLM_R_X15Y131_SLICE_X21Y131_BO6),
.O5(CLBLM_L_X12Y128_SLICE_X16Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X16Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y128_SLICE_X17Y128_AO6),
.Q(CLBLM_L_X12Y128_SLICE_X17Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_DO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_CO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_BO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafafaaaaabafa)
  ) CLBLM_L_X12Y128_SLICE_X17Y128_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_CO6),
.I2(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I3(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_AO6),
.I5(CLBLM_R_X15Y129_SLICE_X21Y129_BQ),
.O5(CLBLM_L_X12Y128_SLICE_X17Y128_AO5),
.O6(CLBLM_L_X12Y128_SLICE_X17Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y129_SLICE_X16Y129_BO6),
.Q(CLBLM_L_X12Y129_SLICE_X16Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77f777f777f7ffff)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_CLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I1(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I2(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I3(CLBLM_R_X15Y129_SLICE_X21Y129_BQ),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555000054545404)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I1(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_CO6),
.I3(CLBLM_L_X12Y129_SLICE_X16Y129_CO6),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_AO6),
.I5(CLBLM_L_X12Y129_SLICE_X16Y129_AO5),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h004000000f4f0f4f)
  ) CLBLM_L_X12Y129_SLICE_X16Y129_ALUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I2(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I4(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X16Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X16Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X18Y129_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y101_IOB_X0Y101_I),
.Q(CLBLM_L_X12Y129_SLICE_X17Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_DO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fcf0f0f0f0f0)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I3(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_CO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaaafaaaeaeafaf)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I1(CLBLM_R_X15Y129_SLICE_X21Y129_BQ),
.I2(CLBLM_L_X12Y129_SLICE_X16Y129_AO6),
.I3(CLBLM_R_X13Y128_SLICE_X18Y128_CO6),
.I4(CLBLM_R_X15Y129_SLICE_X21Y129_DO6),
.I5(CLBLM_L_X12Y129_SLICE_X17Y129_AO5),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_BO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha080a080ffddffff)
  ) CLBLM_L_X12Y129_SLICE_X17Y129_ALUT (
.I0(CLBLM_L_X12Y128_SLICE_X17Y128_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y129_SLICE_X17Y129_AO5),
.O6(CLBLM_L_X12Y129_SLICE_X17Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_AO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_BO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y130_SLICE_X16Y130_CO6),
.Q(CLBLM_L_X12Y130_SLICE_X16Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h11f155f511115555)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_DLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cfc0cfc0cfc0efe)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_CLUT (
.I0(CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR),
.I1(CLBLM_L_X12Y130_SLICE_X17Y130_AO6),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I4(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I5(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f1d3f0c1d1d0c0c)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_BLUT (
.I0(CLBLM_L_X12Y130_SLICE_X16Y130_DO6),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I3(CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_BO6),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444544eeeeefee)
  ) CLBLM_L_X12Y130_SLICE_X16Y130_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I1(CLBLM_L_X10Y130_SLICE_X13Y130_BO6),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I3(CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR),
.I4(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.O5(CLBLM_L_X12Y130_SLICE_X16Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X16Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y101_IOB_X0Y101_I),
.Q(CLBLM_L_X12Y130_SLICE_X17Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_DO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000f0f000000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I5(CLBLM_L_X12Y130_SLICE_X17Y130_BO6),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_CO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000020000000)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_BO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0088000f0f8888)
  ) CLBLM_L_X12Y130_SLICE_X17Y130_ALUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AO6),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_A5Q),
.I4(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I5(CLBLM_L_X12Y130_SLICE_X17Y130_CO6),
.O5(CLBLM_L_X12Y130_SLICE_X17Y130_AO5),
.O6(CLBLM_L_X12Y130_SLICE_X17Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y131_SLICE_X16Y131_AO5),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.Q(CLBLM_L_X12Y131_SLICE_X16Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heaea00eaea400040)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_DLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR),
.I3(CLBLM_L_X12Y130_SLICE_X17Y130_CO6),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_A5Q),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77dd278d72d82288)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_CLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I4(CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cccccccf0000000)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0f0055cc55cc)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_ALUT (
.I0(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_CO6),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y131_SLICE_X17Y131_AO5),
.Q(CLBLM_L_X12Y131_SLICE_X17Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y131_SLICE_X17Y131_AO6),
.Q(CLBLM_L_X12Y131_SLICE_X17Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0005000500050)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_DLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7722777777222222)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_CLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR),
.I4(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0faaccf0f0aacc)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030fcfc22ee22ee)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_ALUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_BO6),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f1b4e0af5b1e4a0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_DLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_L_X12Y132_SLICE_X17Y132_DO6),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_B5Q),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h45efef4540eaea40)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_CLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_AO5),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.I5(CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3022fceefcee3022)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR),
.I1(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_A5Q),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000000080000000)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_A5Q),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y132_SLICE_X17Y132_AO5),
.Q(CLBLM_L_X12Y132_SLICE_X17Y132_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y132_SLICE_X17Y132_BO5),
.Q(CLBLM_L_X12Y132_SLICE_X17Y132_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y132_SLICE_X17Y132_AO6),
.Q(CLBLM_L_X12Y132_SLICE_X17Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y132_SLICE_X17Y132_BO6),
.Q(CLBLM_L_X12Y132_SLICE_X17Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I1(CLBLM_L_X12Y131_SLICE_X17Y131_A5Q),
.I2(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.I3(CLBLM_L_X12Y132_SLICE_X17Y132_A5Q),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h45efef4540eaea40)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_CLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_L_X12Y132_SLICE_X17Y132_A5Q),
.I4(CLBLM_L_X12Y133_SLICE_X17Y133_DO6),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f033f055ff5500)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_BLUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I1(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_CO6),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0dddd8888)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_ALUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.I1(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_CO6),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_BO5),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_AO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_BO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3131f5f531310000)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_DLUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444a0f5a0f5)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I1(CLBLM_R_X13Y133_SLICE_X18Y133_BO5),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_CO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fc00fcccc3ccc3)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_B5Q),
.I2(CLBLM_R_X13Y135_SLICE_X19Y135_DQ),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50f0f0f870f0f0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_ALUT (
.I0(CLBLM_L_X12Y134_SLICE_X16Y134_DO6),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I3(CLBLM_R_X13Y134_SLICE_X18Y134_BO6),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.I5(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.Q(CLBLM_L_X12Y133_SLICE_X17Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888800000000)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3311ff550000cc44)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_CLUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5bbf511a0bba011)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_CO6),
.I5(CLBLM_R_X13Y133_SLICE_X18Y133_BO6),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heecfee0322cf2203)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_ALUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_AO5),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I2(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_CO6),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_CO6),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.Q(CLBLM_L_X12Y134_SLICE_X16Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0ccc00c000c00)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I3(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_BQ),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaa30aa00)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.I2(CLBLM_R_X3Y126_SLICE_X2Y126_AQ),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_CO6),
.I4(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010dfef2ffff)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_BLUT (
.I0(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80808080ff00ff00)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_ALUT (
.I0(CLBLM_L_X12Y134_SLICE_X16Y134_DO6),
.I1(CLBLM_R_X13Y134_SLICE_X18Y134_BO6),
.I2(CLBLM_L_X12Y134_SLICE_X17Y134_CO6),
.I3(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c5c0cfc0cf)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_DLUT (
.I0(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I1(CLBLM_R_X13Y133_SLICE_X18Y133_CO6),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I3(CLBLM_R_X13Y135_SLICE_X19Y135_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000045550111)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I2(CLBLM_R_X3Y126_SLICE_X2Y126_AQ),
.I3(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.I4(CLBLM_R_X15Y137_SLICE_X20Y137_D_CY),
.I5(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8cc00b8b8ff33)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_BO6),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_CO6),
.I3(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I5(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a000000020)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_ALUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_AQ),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I2(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.Q(CLBLM_L_X12Y135_SLICE_X16Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.Q(CLBLM_L_X12Y135_SLICE_X16Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffaf0faf0fa)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_DLUT (
.I0(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_CLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc50ccfacc)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_BLUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3d1f2d0e2c0f2d0)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_ALUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_CO6),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I3(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_CO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_L_X12Y135_SLICE_X17Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00f0cccc0fff)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y135_SLICE_X19Y135_BO6),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I5(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb80000ff000000)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_CLUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_BQ),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.I5(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h474747470033ccff)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_BLUT (
.I0(CLBLM_L_X16Y134_SLICE_X22Y134_AO5),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_AQ),
.I3(CLBLM_L_X12Y137_SLICE_X16Y137_BQ),
.I4(CLBLM_R_X15Y134_SLICE_X20Y134_BQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0dddd8888)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I2(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff3f3000f0303)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y137_SLICE_X18Y137_CO6),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_CO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_BO6),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_DO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ddf588a0dda088)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_CQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_AO5),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.I4(CLBLM_R_X15Y138_SLICE_X21Y138_AQ),
.I5(CLBLM_R_X15Y135_SLICE_X21Y135_AQ),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_CO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccaaaa)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_BLUT (
.I0(CLBLM_R_X15Y137_SLICE_X21Y137_BQ),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_BQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_AO6),
.I3(CLBLM_R_X15Y134_SLICE_X21Y134_CQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_BO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f0f0f00000)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y136_SLICE_X17Y136_AO6),
.Q(CLBLM_L_X12Y136_SLICE_X17Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.Q(CLBLM_L_X12Y136_SLICE_X17Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y136_SLICE_X17Y136_CO6),
.Q(CLBLM_L_X12Y136_SLICE_X17Y136_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1b1b00aa1b1b55ff)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLL_L_X26Y138_SLICE_X38Y138_AO5),
.I3(CLBLM_R_X13Y131_SLICE_X18Y131_DQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.I5(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_DO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ecffec004cff4c)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_CO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffecec4c4c)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_BLUT (
.I0(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.I3(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_BO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fffffc74fc74)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_ALUT (
.I0(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I1(CLBLM_L_X12Y137_SLICE_X17Y137_CO5),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_AO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y137_SLICE_X16Y137_BO6),
.Q(CLBLM_L_X12Y137_SLICE_X16Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f3fffff5f0fffff)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aaaaaa22aa22aa)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_CLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.I2(1'b1),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0cfcccccacac)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X12Y137_SLICE_X16Y137_BQ),
.I2(CLBLM_R_X13Y140_SLICE_X19Y140_AO6),
.I3(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I4(CLBLM_L_X8Y138_SLICE_X11Y138_AO6),
.I5(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055ff5530353f35)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_ALUT (
.I0(CLBLM_R_X13Y138_SLICE_X19Y138_BQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y137_SLICE_X17Y137_AO6),
.Q(CLBLM_L_X12Y137_SLICE_X17Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y137_SLICE_X17Y137_BO6),
.Q(CLBLM_L_X12Y137_SLICE_X17Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_DLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I2(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fff3fffff00aaaa)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_CLUT (
.I0(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.I4(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cacccccfcacccc)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X12Y137_SLICE_X17Y137_BQ),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_CO6),
.I3(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.I4(CLBLM_R_X13Y140_SLICE_X19Y140_AO6),
.I5(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f0f0f0aaf0f0f0)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_AQ),
.I3(CLBLM_R_X13Y140_SLICE_X19Y140_AO6),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_BO6),
.I5(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.DIB(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.DIC(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.DID(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.DOA(CLBLM_L_X12Y138_SLICE_X16Y138_AO6),
.DOB(CLBLM_L_X12Y138_SLICE_X16Y138_BO6),
.DOC(CLBLM_L_X12Y138_SLICE_X16Y138_CO6),
.DOD(CLBLM_L_X12Y138_SLICE_X16Y138_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_R_X11Y139_SLICE_X15Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_CO6),
.Q(CLBLM_L_X12Y138_SLICE_X17Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_DO6),
.Q(CLBLM_L_X12Y138_SLICE_X17Y138_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_DO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_CO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcccccccc)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_BO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddf5dda088f588a0)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_BQ),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I4(CLBLM_L_X12Y137_SLICE_X17Y137_AQ),
.I5(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_AO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X10Y139_SLICE_X13Y139_BO6),
.DIB(CLBLM_R_X13Y142_SLICE_X18Y142_AO6),
.DIC(CLBLM_R_X13Y141_SLICE_X18Y141_CO6),
.DID(1'b0),
.DOA(CLBLM_L_X12Y139_SLICE_X16Y139_AO6),
.DOB(CLBLM_L_X12Y139_SLICE_X16Y139_BO6),
.DOC(CLBLM_L_X12Y139_SLICE_X16Y139_CO6),
.DOD(CLBLM_L_X12Y139_SLICE_X16Y139_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_R_X11Y139_SLICE_X15Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000100010001000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_AO6),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_DO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffe4e4ffff0000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I2(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_CO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaebfffaeaeffff)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_BO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000008000000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_AO6),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_AO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X10Y139_SLICE_X13Y139_BO6),
.DIB(CLBLM_R_X13Y142_SLICE_X18Y142_AO6),
.DIC(CLBLM_R_X13Y141_SLICE_X18Y141_CO6),
.DID(1'b0),
.DOA(CLBLM_L_X12Y140_SLICE_X16Y140_AO6),
.DOB(CLBLM_L_X12Y140_SLICE_X16Y140_BO6),
.DOC(CLBLM_L_X12Y140_SLICE_X16Y140_CO6),
.DOD(CLBLM_L_X12Y140_SLICE_X16Y140_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_L_X12Y140_SLICE_X17Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y140_SLICE_X17Y140_AO6),
.Q(CLBLM_L_X12Y140_SLICE_X17Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y140_SLICE_X17Y140_BO6),
.Q(CLBLM_L_X12Y140_SLICE_X17Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000500000000000)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_AO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_DO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff10ff00ff00)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_CLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_L_X12Y141_SLICE_X17Y141_BO6),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_CO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c0c5500fcacffaa)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_BLUT (
.I0(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_DO6),
.I5(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_BO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccd8ccccccd8d8d8)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_ALUT (
.I0(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_AO6),
.I2(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I3(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_DO6),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_AO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X10Y139_SLICE_X13Y139_BO6),
.DIB(CLBLM_R_X13Y142_SLICE_X18Y142_AO6),
.DIC(CLBLM_R_X13Y141_SLICE_X18Y141_CO6),
.DID(1'b0),
.DOA(CLBLM_L_X12Y141_SLICE_X16Y141_AO6),
.DOB(CLBLM_L_X12Y141_SLICE_X16Y141_BO6),
.DOC(CLBLM_L_X12Y141_SLICE_X16Y141_CO6),
.DOD(CLBLM_L_X12Y141_SLICE_X16Y141_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_L_X12Y139_SLICE_X17Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y141_SLICE_X18Y141_CO6),
.Q(CLBLM_L_X12Y141_SLICE_X17Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f303f3f3030303)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_L_X12Y141_SLICE_X17Y141_AO5),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_CO5),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_DO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5500553f550055)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_CLUT (
.I0(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_CO6),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_CO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888ddd58880)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_AO6),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_BO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a000a00a000a000)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_ALUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_AO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X12Y140_SLICE_X17Y140_CO6),
.DIB(CLBLM_L_X12Y142_SLICE_X17Y142_DO6),
.DIC(CLBLM_R_X13Y141_SLICE_X18Y141_BO6),
.DID(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.DOA(CLBLM_L_X12Y142_SLICE_X16Y142_AO6),
.DOB(CLBLM_L_X12Y142_SLICE_X16Y142_BO6),
.DOC(CLBLM_L_X12Y142_SLICE_X16Y142_CO6),
.DOD(CLBLM_L_X12Y142_SLICE_X16Y142_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_L_X12Y139_SLICE_X17Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_BO5),
.Q(CLBLM_L_X12Y142_SLICE_X17Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y142_SLICE_X17Y142_BO6),
.Q(CLBLM_L_X12Y142_SLICE_X17Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff08ff00)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_DLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I3(CLBLM_L_X12Y142_SLICE_X17Y142_CO6),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_DO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0af808fa0af)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_AO6),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_CO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_BO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00000088880000)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_AO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_AO6),
.Q(CLBLM_L_X12Y143_SLICE_X16Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a0000000)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_DLUT (
.I0(CLBLM_R_X13Y140_SLICE_X19Y140_AO6),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333aaaaf000)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I2(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_CO6),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_DO6),
.I5(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555000000000005)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_BLUT (
.I0(CLBLM_L_X12Y143_SLICE_X16Y143_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff4f4f400b0b0b0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_ALUT (
.I0(CLBLM_L_X12Y137_SLICE_X16Y137_CO5),
.I1(CLBLM_R_X13Y140_SLICE_X19Y140_AO6),
.I2(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.I3(CLBLM_L_X12Y143_SLICE_X16Y143_BO6),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I5(CLBLM_L_X12Y143_SLICE_X16Y143_CO6),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7744444477447474)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_ALUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I1(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.I2(CLBLM_R_X13Y148_SLICE_X18Y148_CO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_DO6),
.I5(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e000e06ff00ff26)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_BO6),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_CO6),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I5(CLBLM_L_X12Y144_SLICE_X16Y144_BO6),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00080808fff7fff7)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacaff0ff000)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_ALUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_B_XOR),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88ff005f0aff00)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_DLUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_AO5),
.I2(CLBLM_R_X13Y145_SLICE_X19Y145_BO5),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a022772277)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_D_XOR),
.I2(CLBLM_R_X13Y144_SLICE_X18Y144_C_XOR),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h114433ecbbee33ec)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb133bb3311331b33)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_L_X12Y144_SLICE_X17Y144_CO5),
.I5(CLBLM_R_X13Y145_SLICE_X19Y145_AO5),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X12Y144_SLICE_X17Y144_MUXF7A (
.I0(CLBLM_L_X12Y144_SLICE_X17Y144_BO6),
.I1(CLBLM_L_X12Y144_SLICE_X17Y144_AO6),
.O(CLBLM_L_X12Y144_SLICE_X17Y144_F7AMUX_O),
.S(CLBLM_R_X15Y150_SLICE_X20Y150_DO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0fff0aaf0ee)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_DLUT (
.I0(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_BO6),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I3(CLBLM_L_X12Y137_SLICE_X17Y137_CO6),
.I4(CLBLM_R_X13Y148_SLICE_X19Y148_BO6),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff8888ffff0a00)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_CLUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I2(CLBLM_L_X10Y148_SLICE_X13Y148_AO5),
.I3(CLBLM_R_X11Y143_SLICE_X15Y143_BO6),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00050c050c050f05)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0000555555ff)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_CO6),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c5fecff4c00eca0)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_DLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_R_X13Y145_SLICE_X18Y145_D_XOR),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0f0e0f0f0f0f)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I2(CLBLM_L_X12Y139_SLICE_X17Y139_BO6),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_BO6),
.I4(CLBLM_R_X13Y148_SLICE_X19Y148_BO6),
.I5(CLBLM_L_X12Y142_SLICE_X17Y142_AO5),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3133313331333131)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_BLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_AO6),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_BO6),
.I2(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I3(CLBLM_R_X13Y148_SLICE_X19Y148_BO6),
.I4(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I5(CLBLM_L_X12Y150_SLICE_X16Y150_BO6),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e00fef00e0efefe)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_ALUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_BO6),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I3(CLBLM_R_X13Y148_SLICE_X19Y148_AO6),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_CO6),
.I5(CLBLM_R_X15Y149_SLICE_X20Y149_CO6),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y152_SLICE_X20Y152_DO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000005500000015)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_DLUT (
.I0(CLBLM_R_X11Y147_SLICE_X15Y147_DO6),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I2(CLBLM_L_X12Y146_SLICE_X17Y146_DO6),
.I3(CLBLM_R_X15Y148_SLICE_X20Y148_AO6),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_DO6),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_BO6),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000acacacac)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_CLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0f000c0c0005)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_BLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafefffffafa)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_DO6),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_DO6),
.I2(CLBLM_R_X15Y148_SLICE_X20Y148_AO6),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_BO6),
.I4(CLBLM_R_X11Y147_SLICE_X15Y147_DO6),
.I5(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fffccff55ff55ff)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_DLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I1(CLBLM_L_X12Y144_SLICE_X17Y144_CO6),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88fcfc3030)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_CLUT (
.I0(CLBLM_L_X12Y144_SLICE_X17Y144_F7AMUX_O),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I2(CLBLM_R_X13Y150_SLICE_X19Y150_F7AMUX_O),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_F7AMUX_O),
.I4(CLBLM_R_X15Y146_SLICE_X21Y146_F7AMUX_O),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020080000000800)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_R_X15Y152_SLICE_X20Y152_DO6),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80a0808000200000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_DO6),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X12Y146_SLICE_X17Y146_MUXF7A (
.I0(CLBLM_L_X12Y146_SLICE_X17Y146_BO6),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_AO6),
.O(CLBLM_L_X12Y146_SLICE_X17Y146_F7AMUX_O),
.S(CLBLM_R_X15Y150_SLICE_X20Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_BQ),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X12Y147_SLICE_X16Y147_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X12Y147_SLICE_X16Y147_D_CY, CLBLM_L_X12Y147_SLICE_X16Y147_C_CY, CLBLM_L_X12Y147_SLICE_X16Y147_B_CY, CLBLM_L_X12Y147_SLICE_X16Y147_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X12Y147_SLICE_X16Y147_DO5, CLBLM_L_X12Y147_SLICE_X16Y147_CO5, CLBLM_L_X12Y147_SLICE_X16Y147_BO5, 1'b0}),
.O({CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR, CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR, CLBLM_L_X12Y147_SLICE_X16Y147_B_XOR, CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR}),
.S({CLBLM_L_X12Y147_SLICE_X16Y147_DO6, CLBLM_L_X12Y147_SLICE_X16Y147_CO6, CLBLM_L_X12Y147_SLICE_X16Y147_BO6, CLBLM_L_X12Y147_SLICE_X16Y147_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h050505fa000000ff)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_DLUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h050505fa000000ff)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_CLUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505363605050505)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f00000f0f)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR),
.Q(CLBLM_L_X12Y147_SLICE_X17Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR),
.Q(CLBLM_L_X12Y147_SLICE_X17Y147_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR),
.Q(CLBLM_L_X12Y147_SLICE_X17Y147_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR),
.Q(CLBLM_L_X12Y147_SLICE_X17Y147_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X12Y147_SLICE_X17Y147_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X12Y147_SLICE_X17Y147_D_CY, CLBLM_L_X12Y147_SLICE_X17Y147_C_CY, CLBLM_L_X12Y147_SLICE_X17Y147_B_CY, CLBLM_L_X12Y147_SLICE_X17Y147_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR, CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR, CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR, 1'b0}),
.O({CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR, CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR, CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR, CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR}),
.S({CLBLM_L_X12Y147_SLICE_X17Y147_DO6, CLBLM_L_X12Y147_SLICE_X17Y147_CO6, CLBLM_L_X12Y147_SLICE_X17Y147_BO6, CLBLM_L_X12Y147_SLICE_X17Y147_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa77887788)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_DLUT (
.I0(CLBLM_L_X12Y147_SLICE_X17Y147_BQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR),
.I4(1'b1),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff0055aaff00)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_CLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR),
.I4(CLBLM_L_X12Y147_SLICE_X17Y147_AQ),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f03c3cf0f0)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR),
.I3(1'b1),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y147_SLICE_X16Y147_B_XOR),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X12Y148_SLICE_X16Y148_CARRY4 (
.CI(CLBLM_L_X12Y147_SLICE_X16Y147_COUT),
.CO({CLBLM_L_X12Y148_SLICE_X16Y148_D_CY, CLBLM_L_X12Y148_SLICE_X16Y148_C_CY, CLBLM_L_X12Y148_SLICE_X16Y148_B_CY, CLBLM_L_X12Y148_SLICE_X16Y148_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X12Y148_SLICE_X16Y148_DO5, CLBLM_L_X12Y148_SLICE_X16Y148_CO5, CLBLM_L_X12Y148_SLICE_X16Y148_BO5, CLBLM_L_X12Y148_SLICE_X16Y148_AO5}),
.O({CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR, CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR, CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR, CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR}),
.S({CLBLM_L_X12Y148_SLICE_X16Y148_DO6, CLBLM_L_X12Y148_SLICE_X16Y148_CO6, CLBLM_L_X12Y148_SLICE_X16Y148_BO6, CLBLM_L_X12Y148_SLICE_X16Y148_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033556600005555)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_DLUT (
.I0(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h111111ee11111111)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_CLUT (
.I0(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033556600005555)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055336600003333)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR),
.Q(CLBLM_L_X12Y148_SLICE_X17Y148_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR),
.Q(CLBLM_L_X12Y148_SLICE_X17Y148_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR),
.Q(CLBLM_L_X12Y148_SLICE_X17Y148_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR),
.Q(CLBLM_L_X12Y148_SLICE_X17Y148_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X12Y148_SLICE_X17Y148_CARRY4 (
.CI(CLBLM_L_X12Y147_SLICE_X17Y147_COUT),
.CO({CLBLM_L_X12Y148_SLICE_X17Y148_D_CY, CLBLM_L_X12Y148_SLICE_X17Y148_C_CY, CLBLM_L_X12Y148_SLICE_X17Y148_B_CY, CLBLM_L_X12Y148_SLICE_X17Y148_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR, CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR, CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR, CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR}),
.O({CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR, CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR, CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR, CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR}),
.S({CLBLM_L_X12Y148_SLICE_X17Y148_DO6, CLBLM_L_X12Y148_SLICE_X17Y148_CO6, CLBLM_L_X12Y148_SLICE_X17Y148_BO6, CLBLM_L_X12Y148_SLICE_X17Y148_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f03f3fc0c0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I2(CLBLM_L_X12Y148_SLICE_X17Y148_BQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa6666aaaa)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_CLUT (
.I0(CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X12Y148_SLICE_X17Y148_AQ),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3cf03cf0)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y147_SLICE_X17Y147_DQ),
.I2(CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc33cccccc)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR),
.I2(1'b1),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I4(CLBLM_L_X12Y147_SLICE_X17Y147_CQ),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X12Y149_SLICE_X16Y149_CARRY4 (
.CI(CLBLM_L_X12Y148_SLICE_X16Y148_COUT),
.CO({CLBLM_L_X12Y149_SLICE_X16Y149_D_CY, CLBLM_L_X12Y149_SLICE_X16Y149_C_CY, CLBLM_L_X12Y149_SLICE_X16Y149_B_CY, CLBLM_L_X12Y149_SLICE_X16Y149_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X12Y149_SLICE_X16Y149_D_XOR, CLBLM_L_X12Y149_SLICE_X16Y149_C_XOR, CLBLM_L_X12Y149_SLICE_X16Y149_B_XOR, CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR}),
.S({CLBLM_L_X12Y149_SLICE_X16Y149_DO6, CLBLM_L_X12Y149_SLICE_X16Y149_CO6, CLBLM_L_X12Y149_SLICE_X16Y149_BO6, CLBLM_L_X12Y149_SLICE_X16Y149_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ff000000ff)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X12Y149_SLICE_X17Y149_CARRY4 (
.CI(CLBLM_L_X12Y148_SLICE_X17Y148_COUT),
.CO({CLBLM_L_X12Y149_SLICE_X17Y149_D_CY, CLBLM_L_X12Y149_SLICE_X17Y149_C_CY, CLBLM_L_X12Y149_SLICE_X17Y149_B_CY, CLBLM_L_X12Y149_SLICE_X17Y149_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, CLBLM_L_X12Y149_SLICE_X16Y149_B_CY}),
.O({CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR, CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR, CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR, CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR}),
.S({CLBLM_L_X12Y149_SLICE_X17Y149_DO6, CLBLM_L_X12Y149_SLICE_X17Y149_CO6, CLBLM_L_X12Y149_SLICE_X17Y149_BO6, CLBLM_L_X12Y149_SLICE_X17Y149_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa88888888)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_DLUT (
.I0(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee0000eeee0000)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_CLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa88888888)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_BLUT (
.I0(CLBLM_L_X12Y148_SLICE_X17Y148_DQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a78787878)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_ALUT (
.I0(CLBLM_L_X12Y148_SLICE_X17Y148_CQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_B_CY),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010001)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_DLUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_DO6),
.I1(CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR),
.I2(CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR),
.I3(CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR),
.I4(1'b1),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f7f557f0a200020)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.I5(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f0f5f1f0f0f0f0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_BLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_AO6),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05055555f00a0f0f)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I3(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR),
.Q(CLBLM_L_X12Y150_SLICE_X17Y150_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X12Y150_SLICE_X17Y150_CARRY4 (
.CI(CLBLM_L_X12Y149_SLICE_X17Y149_COUT),
.CO({CLBLM_L_X12Y150_SLICE_X17Y150_D_CY, CLBLM_L_X12Y150_SLICE_X17Y150_C_CY, CLBLM_L_X12Y150_SLICE_X17Y150_B_CY, CLBLM_L_X12Y150_SLICE_X17Y150_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X12Y150_SLICE_X17Y150_D_XOR, CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR, CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR, CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR}),
.S({CLBLM_L_X12Y150_SLICE_X17Y150_DO6, CLBLM_L_X12Y150_SLICE_X17Y150_CO6, CLBLM_L_X12Y150_SLICE_X17Y150_BO6, CLBLM_L_X12Y150_SLICE_X17Y150_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee0000eeee0000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_CLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaaa0000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_BLUT (
.I0(CLBLM_L_X12Y149_SLICE_X17Y149_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaa00aa00)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_ALUT (
.I0(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a0a0a0a0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5a6a566a565a55)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_CLUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbcf88cfbb038803)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_BLUT (
.I0(CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_AO6),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_CO6),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he1a5f0e1870fa587)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I4(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5fdfdfa0008080)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_DLUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I1(CLBLM_R_X11Y150_SLICE_X15Y150_CO6),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00acac0ff0acac)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_CLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_AO5),
.I1(CLBLM_R_X15Y152_SLICE_X21Y152_CO6),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1b4e33ee1b4e33cc)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h270f270faf0f050f)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_AO6),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X12Y151_SLICE_X17Y151_MUXF7A (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_BO6),
.I1(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.O(CLBLM_L_X12Y151_SLICE_X17Y151_F7AMUX_O),
.S(CLBLM_R_X15Y150_SLICE_X20Y150_DO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X12Y151_SLICE_X17Y151_MUXF7B (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I1(CLBLM_L_X12Y151_SLICE_X17Y151_CO6),
.O(CLBLM_L_X12Y151_SLICE_X17Y151_F7BMUX_O),
.S(CLBLM_R_X15Y150_SLICE_X20Y150_DO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X12Y151_SLICE_X17Y151_MUXF8 (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_F7BMUX_O),
.I1(CLBLM_L_X12Y151_SLICE_X17Y151_F7AMUX_O),
.O(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.S(CLBLM_R_X15Y150_SLICE_X20Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y131_SLICE_X22Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y131_SLICE_X22Y131_AO6),
.Q(CLBLM_L_X16Y131_SLICE_X22Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y131_SLICE_X22Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y131_SLICE_X22Y131_DO5),
.O6(CLBLM_L_X16Y131_SLICE_X22Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y131_SLICE_X22Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y131_SLICE_X22Y131_CO5),
.O6(CLBLM_L_X16Y131_SLICE_X22Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y131_SLICE_X22Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y131_SLICE_X22Y131_BO5),
.O6(CLBLM_L_X16Y131_SLICE_X22Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fcaaaa03ffaaaa)
  ) CLBLM_L_X16Y131_SLICE_X22Y131_ALUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_CQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I3(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I5(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.O5(CLBLM_L_X16Y131_SLICE_X22Y131_AO5),
.O6(CLBLM_L_X16Y131_SLICE_X22Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y131_SLICE_X23Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y131_SLICE_X23Y131_DO5),
.O6(CLBLM_L_X16Y131_SLICE_X23Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y131_SLICE_X23Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y131_SLICE_X23Y131_CO5),
.O6(CLBLM_L_X16Y131_SLICE_X23Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y131_SLICE_X23Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y131_SLICE_X23Y131_BO5),
.O6(CLBLM_L_X16Y131_SLICE_X23Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y131_SLICE_X23Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y131_SLICE_X23Y131_AO5),
.O6(CLBLM_L_X16Y131_SLICE_X23Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y133_SLICE_X22Y133_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y133_SLICE_X22Y133_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y133_SLICE_X22Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y133_SLICE_X22Y133_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y133_SLICE_X22Y133_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y133_SLICE_X22Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y133_SLICE_X22Y133_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y133_SLICE_X22Y133_CO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y133_SLICE_X22Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y133_SLICE_X22Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y133_SLICE_X22Y133_DO5),
.O6(CLBLM_L_X16Y133_SLICE_X22Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0ccf5cccccccc)
  ) CLBLM_L_X16Y133_SLICE_X22Y133_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X16Y133_SLICE_X22Y133_CQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_CO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.O5(CLBLM_L_X16Y133_SLICE_X22Y133_CO5),
.O6(CLBLM_L_X16Y133_SLICE_X22Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaccc0cccacccfcc)
  ) CLBLM_L_X16Y133_SLICE_X22Y133_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X16Y133_SLICE_X22Y133_BQ),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_DO6),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_CO6),
.O5(CLBLM_L_X16Y133_SLICE_X22Y133_BO5),
.O6(CLBLM_L_X16Y133_SLICE_X22Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ddf0f0f011f0)
  ) CLBLM_L_X16Y133_SLICE_X22Y133_ALUT (
.I0(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_L_X16Y133_SLICE_X22Y133_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X16Y133_SLICE_X22Y133_AO5),
.O6(CLBLM_L_X16Y133_SLICE_X22Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y133_SLICE_X23Y133_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y133_SLICE_X23Y133_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y133_SLICE_X23Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y133_SLICE_X23Y133_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y133_SLICE_X23Y133_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y133_SLICE_X23Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y133_SLICE_X23Y133_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y133_SLICE_X23Y133_CO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y133_SLICE_X23Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y133_SLICE_X23Y133_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y133_SLICE_X23Y133_DO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y133_SLICE_X23Y133_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfff37008c0004)
  ) CLBLM_L_X16Y133_SLICE_X23Y133_DLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I3(CLBLM_R_X11Y136_SLICE_X14Y136_DO6),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I5(CLBLM_L_X16Y133_SLICE_X23Y133_DQ),
.O5(CLBLM_L_X16Y133_SLICE_X23Y133_DO5),
.O6(CLBLM_L_X16Y133_SLICE_X23Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000bf378c04)
  ) CLBLM_L_X16Y133_SLICE_X23Y133_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I2(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X16Y133_SLICE_X23Y133_CQ),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_BO6),
.O5(CLBLM_L_X16Y133_SLICE_X23Y133_CO5),
.O6(CLBLM_L_X16Y133_SLICE_X23Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff700c4ff370004)
  ) CLBLM_L_X16Y133_SLICE_X23Y133_BLUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.I4(CLBLM_L_X16Y133_SLICE_X23Y133_BQ),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X16Y133_SLICE_X23Y133_BO5),
.O6(CLBLM_L_X16Y133_SLICE_X23Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4f4b0b0f4b0b0)
  ) CLBLM_L_X16Y133_SLICE_X23Y133_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_CO6),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I2(CLBLM_L_X16Y133_SLICE_X23Y133_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X16Y133_SLICE_X23Y133_AO5),
.O6(CLBLM_L_X16Y133_SLICE_X23Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y134_SLICE_X22Y134_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y134_SLICE_X22Y134_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y134_SLICE_X22Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y134_SLICE_X22Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y134_SLICE_X22Y134_DO5),
.O6(CLBLM_L_X16Y134_SLICE_X22Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccdc8dd88cdc8)
  ) CLBLM_L_X16Y134_SLICE_X22Y134_CLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I1(CLBLM_L_X16Y134_SLICE_X22Y134_AO6),
.I2(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I3(CLBLM_L_X16Y134_SLICE_X22Y134_AO5),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.O5(CLBLM_L_X16Y134_SLICE_X22Y134_CO5),
.O6(CLBLM_L_X16Y134_SLICE_X22Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccd8ccddcc88cc8d)
  ) CLBLM_L_X16Y134_SLICE_X22Y134_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.I1(CLBLM_L_X16Y134_SLICE_X22Y134_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X16Y134_SLICE_X22Y134_BO5),
.O6(CLBLM_L_X16Y134_SLICE_X22Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLM_L_X16Y134_SLICE_X22Y134_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(CLBLM_L_X16Y134_SLICE_X22Y134_BQ),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X16Y135_SLICE_X22Y135_AQ),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(1'b1),
.O5(CLBLM_L_X16Y134_SLICE_X22Y134_AO5),
.O6(CLBLM_L_X16Y134_SLICE_X22Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y134_SLICE_X23Y134_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y134_SLICE_X23Y134_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y134_SLICE_X23Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y134_SLICE_X23Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y134_SLICE_X23Y134_DO5),
.O6(CLBLM_L_X16Y134_SLICE_X23Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y134_SLICE_X23Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y134_SLICE_X23Y134_CO5),
.O6(CLBLM_L_X16Y134_SLICE_X23Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y134_SLICE_X23Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y134_SLICE_X23Y134_BO5),
.O6(CLBLM_L_X16Y134_SLICE_X23Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaf033f0)
  ) CLBLM_L_X16Y134_SLICE_X23Y134_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I2(CLBLM_L_X16Y134_SLICE_X23Y134_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLM_R_X5Y135_SLICE_X6Y135_CO6),
.O5(CLBLM_L_X16Y134_SLICE_X23Y134_AO5),
.O6(CLBLM_L_X16Y134_SLICE_X23Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y135_SLICE_X22Y135_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y135_SLICE_X22Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y135_SLICE_X22Y135_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y135_SLICE_X22Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X22Y135_DO5),
.O6(CLBLM_L_X16Y135_SLICE_X22Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03f3000055550000)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_CLUT (
.I0(CLBLM_L_X16Y136_SLICE_X22Y136_BQ),
.I1(CLBLM_L_X16Y135_SLICE_X22Y135_AQ),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.O5(CLBLM_L_X16Y135_SLICE_X22Y135_CO5),
.O6(CLBLM_L_X16Y135_SLICE_X22Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccca0ccccccaf)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X16Y135_SLICE_X22Y135_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_DO6),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_CO6),
.O5(CLBLM_L_X16Y135_SLICE_X22Y135_BO5),
.O6(CLBLM_L_X16Y135_SLICE_X22Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0bbf088)
  ) CLBLM_L_X16Y135_SLICE_X22Y135_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_L_X16Y135_SLICE_X22Y135_AQ),
.I3(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_CO6),
.O5(CLBLM_L_X16Y135_SLICE_X22Y135_AO5),
.O6(CLBLM_L_X16Y135_SLICE_X22Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y135_SLICE_X23Y135_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y135_SLICE_X23Y135_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y135_SLICE_X23Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y135_SLICE_X23Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X23Y135_DO5),
.O6(CLBLM_L_X16Y135_SLICE_X23Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y135_SLICE_X23Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X23Y135_CO5),
.O6(CLBLM_L_X16Y135_SLICE_X23Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y135_SLICE_X23Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y135_SLICE_X23Y135_BO5),
.O6(CLBLM_L_X16Y135_SLICE_X23Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f0d1f0c0f0d1)
  ) CLBLM_L_X16Y135_SLICE_X23Y135_ALUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.I2(CLBLM_L_X16Y135_SLICE_X23Y135_AQ),
.I3(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X16Y135_SLICE_X23Y135_AO5),
.O6(CLBLM_L_X16Y135_SLICE_X23Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_BO6),
.Q(CLBLM_L_X16Y136_SLICE_X22Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5550555000000000)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y137_SLICE_X19Y137_BQ),
.O5(CLBLM_L_X16Y136_SLICE_X22Y136_DO5),
.O6(CLBLM_L_X16Y136_SLICE_X22Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaaafaaafaaefe)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_CLUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I1(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_CO6),
.I4(CLBLM_L_X16Y136_SLICE_X22Y136_DO6),
.I5(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.O5(CLBLM_L_X16Y136_SLICE_X22Y136_CO5),
.O6(CLBLM_L_X16Y136_SLICE_X22Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff50f05cccccccc)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_BLUT (
.I0(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I1(CLBLM_L_X16Y136_SLICE_X22Y136_BQ),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I5(CLBLM_L_X16Y136_SLICE_X22Y136_CO6),
.O5(CLBLM_L_X16Y136_SLICE_X22Y136_BO5),
.O6(CLBLM_L_X16Y136_SLICE_X22Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0fdd88)
  ) CLBLM_L_X16Y136_SLICE_X22Y136_ALUT (
.I0(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I3(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y136_SLICE_X22Y136_AO5),
.O6(CLBLM_L_X16Y136_SLICE_X22Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X23Y136_AO6),
.Q(CLBLM_L_X16Y136_SLICE_X23Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y136_SLICE_X23Y136_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y136_SLICE_X23Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y136_SLICE_X23Y136_CO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y136_SLICE_X23Y136_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y136_SLICE_X23Y136_DO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y136_SLICE_X23Y136_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b8f0fcf030f074)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_DLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.I2(CLBLM_L_X16Y136_SLICE_X23Y136_DQ),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X16Y136_SLICE_X23Y136_DO5),
.O6(CLBLM_L_X16Y136_SLICE_X23Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccccf5cc05)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_CLUT (
.I0(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I1(CLBLM_L_X16Y136_SLICE_X23Y136_CQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_CO6),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I5(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.O5(CLBLM_L_X16Y136_SLICE_X23Y136_CO5),
.O6(CLBLM_L_X16Y136_SLICE_X23Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefcfffd02000301)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_BO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I5(CLBLM_L_X16Y136_SLICE_X23Y136_BQ),
.O5(CLBLM_L_X16Y136_SLICE_X23Y136_BO5),
.O6(CLBLM_L_X16Y136_SLICE_X23Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0f0f0)
  ) CLBLM_L_X16Y136_SLICE_X23Y136_ALUT (
.I0(CLBLM_L_X16Y136_SLICE_X22Y136_AO5),
.I1(1'b1),
.I2(CLBLM_L_X16Y136_SLICE_X23Y136_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X13Y136_SLICE_X19Y136_DO6),
.O5(CLBLM_L_X16Y136_SLICE_X23Y136_AO5),
.O6(CLBLM_L_X16Y136_SLICE_X23Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff084cfdec)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_DLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_L_X16Y137_SLICE_X23Y137_AO6),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I4(CLBLM_L_X16Y137_SLICE_X22Y137_BO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_L_X16Y137_SLICE_X22Y137_DO5),
.O6(CLBLM_L_X16Y137_SLICE_X22Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaacacaacc)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_CLUT (
.I0(CLBLM_L_X16Y137_SLICE_X22Y137_AO6),
.I1(CLBLL_L_X26Y136_SLICE_X38Y136_AO5),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_L_X16Y137_SLICE_X22Y137_CO5),
.O6(CLBLM_L_X16Y137_SLICE_X22Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0fdec3120)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(RIOB33_X105Y119_IOB_X1Y120_I),
.I3(CLBLM_L_X16Y138_SLICE_X22Y138_AQ),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X22Y137_BO5),
.O6(CLBLM_L_X16Y137_SLICE_X22Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22227777f0ddf088)
  ) CLBLM_L_X16Y137_SLICE_X22Y137_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(RIOB33_X105Y121_IOB_X1Y122_I),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I4(CLBLM_L_X16Y137_SLICE_X23Y137_CQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X22Y137_AO5),
.O6(CLBLM_L_X16Y137_SLICE_X22Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y137_SLICE_X23Y137_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y137_SLICE_X23Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y137_SLICE_X23Y137_CO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y137_SLICE_X23Y137_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X23Y137_DO5),
.O6(CLBLM_L_X16Y137_SLICE_X23Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccce4eecccc444e)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_CLUT (
.I0(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.I1(CLBLM_L_X16Y137_SLICE_X23Y137_CQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_DO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X16Y137_SLICE_X23Y137_CO5),
.O6(CLBLM_L_X16Y137_SLICE_X23Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccac0cfc5c)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X16Y137_SLICE_X23Y137_BQ),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I5(CLBLM_R_X5Y135_SLICE_X6Y135_CO6),
.O5(CLBLM_L_X16Y137_SLICE_X23Y137_BO5),
.O6(CLBLM_L_X16Y137_SLICE_X23Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111bbbb0f110fbb)
  ) CLBLM_L_X16Y137_SLICE_X23Y137_ALUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I1(CLBLM_L_X16Y137_SLICE_X23Y137_BQ),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X16Y137_SLICE_X23Y137_AO5),
.O6(CLBLM_L_X16Y137_SLICE_X23Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y138_SLICE_X22Y138_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y138_SLICE_X22Y138_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y138_SLICE_X22Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y138_SLICE_X22Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y138_SLICE_X22Y138_DO5),
.O6(CLBLM_L_X16Y138_SLICE_X22Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y138_SLICE_X22Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y138_SLICE_X22Y138_CO5),
.O6(CLBLM_L_X16Y138_SLICE_X22Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y138_SLICE_X22Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y138_SLICE_X22Y138_BO5),
.O6(CLBLM_L_X16Y138_SLICE_X22Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0bbf0f0f011f0f0)
  ) CLBLM_L_X16Y138_SLICE_X22Y138_ALUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I2(CLBLM_L_X16Y138_SLICE_X22Y138_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_BO6),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_L_X16Y138_SLICE_X22Y138_AO5),
.O6(CLBLM_L_X16Y138_SLICE_X22Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y138_SLICE_X23Y138_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y138_SLICE_X23Y138_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y138_SLICE_X23Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y138_SLICE_X23Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y138_SLICE_X23Y138_DO5),
.O6(CLBLM_L_X16Y138_SLICE_X23Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y138_SLICE_X23Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y138_SLICE_X23Y138_CO5),
.O6(CLBLM_L_X16Y138_SLICE_X23Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y138_SLICE_X23Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y138_SLICE_X23Y138_BO5),
.O6(CLBLM_L_X16Y138_SLICE_X23Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f088f0f0f0dd)
  ) CLBLM_L_X16Y138_SLICE_X23Y138_ALUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_L_X16Y138_SLICE_X23Y138_AQ),
.I3(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_DO6),
.I5(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.O5(CLBLM_L_X16Y138_SLICE_X23Y138_AO5),
.O6(CLBLM_L_X16Y138_SLICE_X23Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y139_SLICE_X22Y139_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y139_SLICE_X22Y139_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y139_SLICE_X22Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y139_SLICE_X22Y139_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X16Y139_SLICE_X22Y139_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_L_X16Y139_SLICE_X22Y139_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y139_SLICE_X22Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y139_SLICE_X22Y139_DO5),
.O6(CLBLM_L_X16Y139_SLICE_X22Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y139_SLICE_X22Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y139_SLICE_X22Y139_CO5),
.O6(CLBLM_L_X16Y139_SLICE_X22Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccac0cfc5c)
  ) CLBLM_L_X16Y139_SLICE_X22Y139_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X16Y139_SLICE_X22Y139_BQ),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_CO6),
.O5(CLBLM_L_X16Y139_SLICE_X22Y139_BO5),
.O6(CLBLM_L_X16Y139_SLICE_X22Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0bbf011)
  ) CLBLM_L_X16Y139_SLICE_X22Y139_ALUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I2(CLBLM_L_X16Y139_SLICE_X22Y139_AQ),
.I3(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_CO6),
.O5(CLBLM_L_X16Y139_SLICE_X22Y139_AO5),
.O6(CLBLM_L_X16Y139_SLICE_X22Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y139_SLICE_X23Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y139_SLICE_X23Y139_DO5),
.O6(CLBLM_L_X16Y139_SLICE_X23Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y139_SLICE_X23Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y139_SLICE_X23Y139_CO5),
.O6(CLBLM_L_X16Y139_SLICE_X23Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y139_SLICE_X23Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y139_SLICE_X23Y139_BO5),
.O6(CLBLM_L_X16Y139_SLICE_X23Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y139_SLICE_X23Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y139_SLICE_X23Y139_AO5),
.O6(CLBLM_L_X16Y139_SLICE_X23Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y140_SLICE_X22Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y143_SLICE_X22Y143_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_L_X16Y140_SLICE_X22Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y140_SLICE_X22Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y143_SLICE_X22Y143_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_L_X16Y140_SLICE_X22Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y140_SLICE_X22Y140_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y143_SLICE_X22Y143_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_L_X16Y140_SLICE_X22Y140_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y140_SLICE_X22Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y140_SLICE_X22Y140_DO5),
.O6(CLBLM_L_X16Y140_SLICE_X22Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y140_SLICE_X22Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y140_SLICE_X22Y140_CO5),
.O6(CLBLM_L_X16Y140_SLICE_X22Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y140_SLICE_X22Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y140_SLICE_X22Y140_BO5),
.O6(CLBLM_L_X16Y140_SLICE_X22Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y140_SLICE_X22Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y140_SLICE_X22Y140_AO5),
.O6(CLBLM_L_X16Y140_SLICE_X22Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y140_SLICE_X23Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y140_SLICE_X23Y140_DO5),
.O6(CLBLM_L_X16Y140_SLICE_X23Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y140_SLICE_X23Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y140_SLICE_X23Y140_CO5),
.O6(CLBLM_L_X16Y140_SLICE_X23Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y140_SLICE_X23Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y140_SLICE_X23Y140_BO5),
.O6(CLBLM_L_X16Y140_SLICE_X23Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y140_SLICE_X23Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y140_SLICE_X23Y140_AO5),
.O6(CLBLM_L_X16Y140_SLICE_X23Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y141_SLICE_X22Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_L_X16Y141_SLICE_X22Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y141_SLICE_X22Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_L_X16Y141_SLICE_X22Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y141_SLICE_X22Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_L_X16Y141_SLICE_X22Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y141_SLICE_X22Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y141_SLICE_X22Y141_DO5),
.O6(CLBLM_L_X16Y141_SLICE_X22Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h030503f5f305f3f5)
  ) CLBLM_L_X16Y141_SLICE_X22Y141_CLUT (
.I0(CLBLM_R_X15Y141_SLICE_X20Y141_CQ),
.I1(CLBLM_L_X16Y141_SLICE_X22Y141_AQ),
.I2(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X15Y141_SLICE_X21Y141_CQ),
.I5(CLBLM_L_X16Y141_SLICE_X23Y141_BQ),
.O5(CLBLM_L_X16Y141_SLICE_X22Y141_CO5),
.O6(CLBLM_L_X16Y141_SLICE_X22Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000000000)
  ) CLBLM_L_X16Y141_SLICE_X22Y141_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_L_X16Y141_SLICE_X22Y141_BO5),
.O6(CLBLM_L_X16Y141_SLICE_X22Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000000)
  ) CLBLM_L_X16Y141_SLICE_X22Y141_ALUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I5(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.O5(CLBLM_L_X16Y141_SLICE_X22Y141_AO5),
.O6(CLBLM_L_X16Y141_SLICE_X22Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y141_SLICE_X23Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y142_SLICE_X22Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_L_X16Y141_SLICE_X23Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y141_SLICE_X23Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y142_SLICE_X22Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_L_X16Y141_SLICE_X23Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y141_SLICE_X23Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y142_SLICE_X22Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_L_X16Y141_SLICE_X23Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y141_SLICE_X23Y141_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y142_SLICE_X22Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_L_X16Y141_SLICE_X23Y141_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y141_SLICE_X23Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y141_SLICE_X23Y141_DO5),
.O6(CLBLM_L_X16Y141_SLICE_X23Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y141_SLICE_X23Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y141_SLICE_X23Y141_CO5),
.O6(CLBLM_L_X16Y141_SLICE_X23Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y141_SLICE_X23Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y141_SLICE_X23Y141_BO5),
.O6(CLBLM_L_X16Y141_SLICE_X23Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y141_SLICE_X23Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y141_SLICE_X23Y141_AO5),
.O6(CLBLM_L_X16Y141_SLICE_X23Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y142_SLICE_X22Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y142_SLICE_X22Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.Q(CLBLM_L_X16Y142_SLICE_X22Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y142_SLICE_X22Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y142_SLICE_X22Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.Q(CLBLM_L_X16Y142_SLICE_X22Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y142_SLICE_X22Y142_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y142_SLICE_X22Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.Q(CLBLM_L_X16Y142_SLICE_X22Y142_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y142_SLICE_X22Y142_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y142_SLICE_X22Y142_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_L_X16Y142_SLICE_X22Y142_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c113f110cdd3fdd)
  ) CLBLM_L_X16Y142_SLICE_X22Y142_DLUT (
.I0(CLBLM_L_X16Y142_SLICE_X23Y142_AQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLM_L_X16Y142_SLICE_X22Y142_AQ),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_AQ),
.I5(CLBLM_R_X15Y142_SLICE_X21Y142_AQ),
.O5(CLBLM_L_X16Y142_SLICE_X22Y142_DO5),
.O6(CLBLM_L_X16Y142_SLICE_X22Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLM_L_X16Y142_SLICE_X22Y142_CLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_L_X16Y142_SLICE_X22Y142_CO5),
.O6(CLBLM_L_X16Y142_SLICE_X22Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c000f3008800bb)
  ) CLBLM_L_X16Y142_SLICE_X22Y142_BLUT (
.I0(CLBLM_R_X15Y144_SLICE_X21Y144_AQ),
.I1(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I2(CLBLM_L_X16Y142_SLICE_X22Y142_AQ),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I4(CLBLM_L_X16Y142_SLICE_X22Y142_AO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_L_X16Y142_SLICE_X22Y142_BO5),
.O6(CLBLM_L_X16Y142_SLICE_X22Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f00fffc0c0c0c0)
  ) CLBLM_L_X16Y142_SLICE_X22Y142_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLM_R_X15Y142_SLICE_X21Y142_AQ),
.I4(CLBLM_L_X16Y142_SLICE_X23Y142_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y142_SLICE_X22Y142_AO5),
.O6(CLBLM_L_X16Y142_SLICE_X22Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y142_SLICE_X23Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.Q(CLBLM_L_X16Y142_SLICE_X23Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y142_SLICE_X23Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y142_SLICE_X23Y142_DO5),
.O6(CLBLM_L_X16Y142_SLICE_X23Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y142_SLICE_X23Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y142_SLICE_X23Y142_CO5),
.O6(CLBLM_L_X16Y142_SLICE_X23Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y142_SLICE_X23Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y142_SLICE_X23Y142_BO5),
.O6(CLBLM_L_X16Y142_SLICE_X23Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y142_SLICE_X23Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y142_SLICE_X23Y142_AO5),
.O6(CLBLM_L_X16Y142_SLICE_X23Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y143_SLICE_X22Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y143_SLICE_X22Y143_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.Q(CLBLM_L_X16Y143_SLICE_X22Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y143_SLICE_X22Y143_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y143_SLICE_X22Y143_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_L_X16Y143_SLICE_X22Y143_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y143_SLICE_X22Y143_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y143_SLICE_X22Y143_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_L_X16Y143_SLICE_X22Y143_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y143_SLICE_X22Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y143_SLICE_X22Y143_DO5),
.O6(CLBLM_L_X16Y143_SLICE_X22Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y143_SLICE_X22Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y143_SLICE_X22Y143_CO5),
.O6(CLBLM_L_X16Y143_SLICE_X22Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y143_SLICE_X22Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y143_SLICE_X22Y143_BO5),
.O6(CLBLM_L_X16Y143_SLICE_X22Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000000000)
  ) CLBLM_L_X16Y143_SLICE_X22Y143_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.O5(CLBLM_L_X16Y143_SLICE_X22Y143_AO5),
.O6(CLBLM_L_X16Y143_SLICE_X22Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y143_SLICE_X23Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y143_SLICE_X23Y143_DO5),
.O6(CLBLM_L_X16Y143_SLICE_X23Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y143_SLICE_X23Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y143_SLICE_X23Y143_CO5),
.O6(CLBLM_L_X16Y143_SLICE_X23Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y143_SLICE_X23Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y143_SLICE_X23Y143_BO5),
.O6(CLBLM_L_X16Y143_SLICE_X23Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y143_SLICE_X23Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y143_SLICE_X23Y143_AO5),
.O6(CLBLM_L_X16Y143_SLICE_X23Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X16Y150_SLICE_X22Y150_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X16Y150_SLICE_X22Y150_D_CY, CLBLM_L_X16Y150_SLICE_X22Y150_C_CY, CLBLM_L_X16Y150_SLICE_X22Y150_B_CY, CLBLM_L_X16Y150_SLICE_X22Y150_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_L_X16Y150_SLICE_X23Y150_CO6, CLBLM_R_X15Y150_SLICE_X21Y150_DO6, CLBLM_L_X16Y150_SLICE_X23Y150_DO6, 1'b0}),
.O({CLBLM_L_X16Y150_SLICE_X22Y150_D_XOR, CLBLM_L_X16Y150_SLICE_X22Y150_C_XOR, CLBLM_L_X16Y150_SLICE_X22Y150_B_XOR, CLBLM_L_X16Y150_SLICE_X22Y150_A_XOR}),
.S({CLBLM_L_X16Y150_SLICE_X22Y150_DO6, CLBLM_L_X16Y150_SLICE_X22Y150_CO6, CLBLM_L_X16Y150_SLICE_X22Y150_BO6, CLBLM_L_X16Y150_SLICE_X22Y150_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc33cc369c33c96)
  ) CLBLM_L_X16Y150_SLICE_X22Y150_DLUT (
.I0(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I1(CLBLM_L_X16Y150_SLICE_X23Y150_CO6),
.I2(CLBLM_L_X16Y150_SLICE_X23Y150_BO5),
.I3(CLBLM_R_X15Y152_SLICE_X21Y152_BQ),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I5(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.O5(CLBLM_L_X16Y150_SLICE_X22Y150_DO5),
.O6(CLBLM_L_X16Y150_SLICE_X22Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc33cc369c33c96)
  ) CLBLM_L_X16Y150_SLICE_X22Y150_CLUT (
.I0(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I1(CLBLM_L_X16Y150_SLICE_X23Y150_AO5),
.I2(CLBLM_R_X15Y150_SLICE_X21Y150_DO6),
.I3(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I5(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.O5(CLBLM_L_X16Y150_SLICE_X22Y150_CO5),
.O6(CLBLM_L_X16Y150_SLICE_X22Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc333cc3c636c636)
  ) CLBLM_L_X16Y150_SLICE_X22Y150_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I1(CLBLM_L_X16Y150_SLICE_X23Y150_DO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_A5Q),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_L_X16Y150_SLICE_X22Y150_BO5),
.O6(CLBLM_L_X16Y150_SLICE_X22Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5f0a5f0f000f0ff)
  ) CLBLM_L_X16Y150_SLICE_X22Y150_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I1(1'b1),
.I2(CLBLM_R_X15Y152_SLICE_X21Y152_AQ),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_L_X16Y150_SLICE_X22Y150_AO5),
.O6(CLBLM_L_X16Y150_SLICE_X22Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafffffffaffffff)
  ) CLBLM_L_X16Y150_SLICE_X23Y150_DLUT (
.I0(CLBLM_R_X15Y152_SLICE_X21Y152_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y150_SLICE_X23Y150_DO5),
.O6(CLBLM_L_X16Y150_SLICE_X23Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf500a000bb11bb11)
  ) CLBLM_L_X16Y150_SLICE_X23Y150_CLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I3(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_L_X16Y150_SLICE_X23Y150_CO5),
.O6(CLBLM_L_X16Y150_SLICE_X23Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfd58f850050a0f0)
  ) CLBLM_L_X16Y150_SLICE_X23Y150_BLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I5(1'b1),
.O5(CLBLM_L_X16Y150_SLICE_X23Y150_BO5),
.O6(CLBLM_L_X16Y150_SLICE_X23Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccaaff55003300)
  ) CLBLM_L_X16Y150_SLICE_X23Y150_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y150_SLICE_X23Y150_AO5),
.O6(CLBLM_L_X16Y150_SLICE_X23Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X16Y151_SLICE_X22Y151_CARRY4 (
.CI(CLBLM_L_X16Y150_SLICE_X22Y150_COUT),
.CO({CLBLM_L_X16Y151_SLICE_X22Y151_D_CY, CLBLM_L_X16Y151_SLICE_X22Y151_C_CY, CLBLM_L_X16Y151_SLICE_X22Y151_B_CY, CLBLM_L_X16Y151_SLICE_X22Y151_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, CLBLM_L_X16Y151_SLICE_X23Y151_BO6, CLBLM_L_X16Y151_SLICE_X23Y151_CO6, CLBLM_L_X16Y151_SLICE_X23Y151_AO6}),
.O({CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR, CLBLM_L_X16Y151_SLICE_X22Y151_C_XOR, CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR, CLBLM_L_X16Y151_SLICE_X22Y151_A_XOR}),
.S({CLBLM_L_X16Y151_SLICE_X22Y151_DO6, CLBLM_L_X16Y151_SLICE_X22Y151_CO6, CLBLM_L_X16Y151_SLICE_X22Y151_BO6, CLBLM_L_X16Y151_SLICE_X22Y151_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f3fff3f0f)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y151_SLICE_X20Y151_BQ),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_CO6),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_L_X16Y151_SLICE_X22Y151_DO5),
.O6(CLBLM_L_X16Y151_SLICE_X22Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c33c3cc3663c99)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_CLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I1(CLBLM_L_X16Y151_SLICE_X23Y151_BO6),
.I2(CLBLM_R_X15Y151_SLICE_X20Y151_BQ),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I4(CLBLM_R_X15Y151_SLICE_X21Y151_CO6),
.I5(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.O5(CLBLM_L_X16Y151_SLICE_X22Y151_CO5),
.O6(CLBLM_L_X16Y151_SLICE_X22Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3963c3cc3c33c69)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_BLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_L_X16Y150_SLICE_X23Y150_BO6),
.I2(CLBLM_L_X16Y151_SLICE_X23Y151_CO6),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I4(CLBLM_L_X16Y151_SLICE_X23Y151_AQ),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.O5(CLBLM_L_X16Y151_SLICE_X22Y151_BO5),
.O6(CLBLM_L_X16Y151_SLICE_X22Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a55a5aa53c5ac3)
  ) CLBLM_L_X16Y151_SLICE_X22Y151_ALUT (
.I0(CLBLM_R_X15Y152_SLICE_X20Y152_AQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I2(CLBLM_L_X16Y151_SLICE_X23Y151_AO6),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I4(CLBLM_L_X16Y150_SLICE_X23Y150_AO6),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_L_X16Y151_SLICE_X22Y151_AO5),
.O6(CLBLM_L_X16Y151_SLICE_X22Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y152_SLICE_X23Y152_BO6),
.Q(CLBLM_L_X16Y151_SLICE_X23Y151_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y151_SLICE_X23Y151_DO5),
.O6(CLBLM_L_X16Y151_SLICE_X23Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8a80000aaaa0202)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_CLUT (
.I0(CLBLM_L_X16Y150_SLICE_X23Y150_AO6),
.I1(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I3(1'b1),
.I4(CLBLM_R_X15Y152_SLICE_X20Y152_AQ),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.O5(CLBLM_L_X16Y151_SLICE_X23Y151_CO5),
.O6(CLBLM_L_X16Y151_SLICE_X23Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000b100b100)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_BLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I2(CLBLM_L_X16Y151_SLICE_X23Y151_AQ),
.I3(CLBLM_L_X16Y150_SLICE_X23Y150_BO6),
.I4(1'b1),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_L_X16Y151_SLICE_X23Y151_BO5),
.O6(CLBLM_L_X16Y151_SLICE_X23Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd008800af05af05)
  ) CLBLM_L_X16Y151_SLICE_X23Y151_ALUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(CLBLM_R_X15Y152_SLICE_X21Y152_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_L_X16Y151_SLICE_X23Y151_AO5),
.O6(CLBLM_L_X16Y151_SLICE_X23Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X16Y152_SLICE_X22Y152_CARRY4 (
.CI(1'b0),
.CO({CLBLM_L_X16Y152_SLICE_X22Y152_D_CY, CLBLM_L_X16Y152_SLICE_X22Y152_C_CY, CLBLM_L_X16Y152_SLICE_X22Y152_B_CY, CLBLM_L_X16Y152_SLICE_X22Y152_A_CY}),
.CYINIT(1'b1),
.DI({CLBLM_R_X15Y150_SLICE_X21Y150_CO6, CLBLM_R_X15Y152_SLICE_X21Y152_AO6, CLBLM_L_X16Y152_SLICE_X23Y152_DO6, CLBLM_L_X16Y152_SLICE_X22Y152_AO5}),
.O({CLBLM_L_X16Y152_SLICE_X22Y152_D_XOR, CLBLM_L_X16Y152_SLICE_X22Y152_C_XOR, CLBLM_L_X16Y152_SLICE_X22Y152_B_XOR, CLBLM_L_X16Y152_SLICE_X22Y152_A_XOR}),
.S({CLBLM_L_X16Y152_SLICE_X22Y152_DO6, CLBLM_L_X16Y152_SLICE_X22Y152_CO6, CLBLM_L_X16Y152_SLICE_X22Y152_BO6, CLBLM_L_X16Y152_SLICE_X22Y152_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h565556559a559a55)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_DLUT (
.I0(CLBLM_R_X15Y150_SLICE_X21Y150_CO6),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_DO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0dd0f22f0110fee)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I1(CLBLM_R_X15Y153_SLICE_X21Y153_AO6),
.I2(CLBLM_L_X16Y150_SLICE_X22Y150_B_XOR),
.I3(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I4(CLBLM_L_X16Y150_SLICE_X23Y150_AO5),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_A5Q),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_CO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f878700ff8877)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_BLUT (
.I0(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I2(CLBLM_L_X16Y150_SLICE_X22Y150_A_XOR),
.I3(CLBLM_R_X15Y152_SLICE_X21Y152_DO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I5(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_BO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1908f7e6eeff0011)
  ) CLBLM_L_X16Y152_SLICE_X22Y152_ALUT (
.I0(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I4(CLBLM_L_X16Y152_SLICE_X23Y152_AQ),
.I5(1'b1),
.O5(CLBLM_L_X16Y152_SLICE_X22Y152_AO5),
.O6(CLBLM_L_X16Y152_SLICE_X22Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y152_SLICE_X23Y152_AO6),
.Q(CLBLM_L_X16Y152_SLICE_X23Y152_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceccceccc4ccc4c)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_DLUT (
.I0(CLBLM_R_X15Y151_SLICE_X20Y151_DO6),
.I1(CLBLM_R_X15Y152_SLICE_X21Y152_DO6),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_DO6),
.I3(CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR),
.I4(1'b1),
.I5(CLBLM_L_X16Y150_SLICE_X22Y150_A_XOR),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_DO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfffdf00800080)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_CLUT (
.I0(CLBLM_R_X15Y151_SLICE_X20Y151_DO6),
.I1(CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_DO6),
.I3(CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR),
.I4(1'b1),
.I5(CLBLM_L_X16Y153_SLICE_X23Y153_BO6),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_CO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0ff00e4e4ff00)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_BLUT (
.I0(CLBLM_L_X16Y154_SLICE_X22Y154_A_CY),
.I1(CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR),
.I2(CLBLM_L_X16Y153_SLICE_X22Y153_C_XOR),
.I3(CLBLM_L_X16Y153_SLICE_X23Y153_BO6),
.I4(CLBLM_R_X15Y151_SLICE_X20Y151_DO6),
.I5(CLBLM_L_X16Y153_SLICE_X23Y153_AO5),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_BO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8b8b888bb)
  ) CLBLM_L_X16Y152_SLICE_X23Y152_ALUT (
.I0(CLBLM_L_X16Y152_SLICE_X22Y152_A_XOR),
.I1(CLBLM_R_X15Y152_SLICE_X20Y152_DO6),
.I2(CLBLM_L_X16Y152_SLICE_X23Y152_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_L_X16Y152_SLICE_X23Y152_AO5),
.O6(CLBLM_L_X16Y152_SLICE_X23Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X16Y153_SLICE_X22Y153_CARRY4 (
.CI(CLBLM_L_X16Y152_SLICE_X22Y152_COUT),
.CO({CLBLM_L_X16Y153_SLICE_X22Y153_D_CY, CLBLM_L_X16Y153_SLICE_X22Y153_C_CY, CLBLM_L_X16Y153_SLICE_X22Y153_B_CY, CLBLM_L_X16Y153_SLICE_X22Y153_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X15Y151_SLICE_X21Y151_BO6, CLBLM_L_X16Y152_SLICE_X23Y152_CO6, CLBLM_R_X15Y152_SLICE_X20Y152_AO6, CLBLM_R_X15Y153_SLICE_X21Y153_BO6}),
.O({CLBLM_L_X16Y153_SLICE_X22Y153_D_XOR, CLBLM_L_X16Y153_SLICE_X22Y153_C_XOR, CLBLM_L_X16Y153_SLICE_X22Y153_B_XOR, CLBLM_L_X16Y153_SLICE_X22Y153_A_XOR}),
.S({CLBLM_L_X16Y153_SLICE_X22Y153_DO6, CLBLM_L_X16Y153_SLICE_X22Y153_CO6, CLBLM_L_X16Y153_SLICE_X22Y153_BO6, CLBLM_L_X16Y153_SLICE_X22Y153_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_L_X16Y153_SLICE_X22Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_BO6),
.O5(CLBLM_L_X16Y153_SLICE_X22Y153_DO5),
.O6(CLBLM_L_X16Y153_SLICE_X22Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d1de2e23f0cc0f3)
  ) CLBLM_L_X16Y153_SLICE_X22Y153_CLUT (
.I0(CLBLM_L_X16Y151_SLICE_X23Y151_AQ),
.I1(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I2(CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I4(CLBLM_R_X15Y151_SLICE_X21Y151_CO6),
.I5(CLBLM_R_X15Y153_SLICE_X21Y153_AO6),
.O5(CLBLM_L_X16Y153_SLICE_X22Y153_CO5),
.O6(CLBLM_L_X16Y153_SLICE_X22Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h028afd7546ceb931)
  ) CLBLM_L_X16Y153_SLICE_X22Y153_BLUT (
.I0(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I4(CLBLM_R_X15Y152_SLICE_X20Y152_AO6),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.O5(CLBLM_L_X16Y153_SLICE_X22Y153_BO5),
.O6(CLBLM_L_X16Y153_SLICE_X22Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03f3fc0c0afaf505)
  ) CLBLM_L_X16Y153_SLICE_X22Y153_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I1(CLBLM_R_X15Y152_SLICE_X21Y152_BQ),
.I2(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I3(CLBLM_L_X16Y150_SLICE_X22Y150_D_XOR),
.I4(CLBLM_L_X16Y150_SLICE_X23Y150_AO6),
.I5(CLBLM_R_X15Y153_SLICE_X21Y153_AO6),
.O5(CLBLM_L_X16Y153_SLICE_X22Y153_AO5),
.O6(CLBLM_L_X16Y153_SLICE_X22Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X23Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X23Y153_DO5),
.O6(CLBLM_L_X16Y153_SLICE_X23Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y153_SLICE_X23Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X23Y153_CO5),
.O6(CLBLM_L_X16Y153_SLICE_X23Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f000f0f0f0ff)
  ) CLBLM_L_X16Y153_SLICE_X23Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X16Y151_SLICE_X23Y151_AQ),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.O5(CLBLM_L_X16Y153_SLICE_X23Y153_BO5),
.O6(CLBLM_L_X16Y153_SLICE_X23Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h20202020dddddddd)
  ) CLBLM_L_X16Y153_SLICE_X23Y153_ALUT (
.I0(CLBLM_R_X15Y151_SLICE_X21Y151_DO6),
.I1(CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR),
.I2(CLBLM_R_X15Y151_SLICE_X20Y151_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y153_SLICE_X23Y153_AO5),
.O6(CLBLM_L_X16Y153_SLICE_X23Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_L_X16Y154_SLICE_X22Y154_CARRY4 (
.CI(CLBLM_L_X16Y153_SLICE_X22Y153_COUT),
.CO({CLBLM_L_X16Y154_SLICE_X22Y154_D_CY, CLBLM_L_X16Y154_SLICE_X22Y154_C_CY, CLBLM_L_X16Y154_SLICE_X22Y154_B_CY, CLBLM_L_X16Y154_SLICE_X22Y154_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_L_X16Y154_SLICE_X22Y154_D_XOR, CLBLM_L_X16Y154_SLICE_X22Y154_C_XOR, CLBLM_L_X16Y154_SLICE_X22Y154_B_XOR, CLBLM_L_X16Y154_SLICE_X22Y154_A_XOR}),
.S({CLBLM_L_X16Y154_SLICE_X22Y154_DO6, CLBLM_L_X16Y154_SLICE_X22Y154_CO6, CLBLM_L_X16Y154_SLICE_X22Y154_BO6, CLBLM_L_X16Y154_SLICE_X22Y154_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X22Y154_DO5),
.O6(CLBLM_L_X16Y154_SLICE_X22Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X22Y154_CO5),
.O6(CLBLM_L_X16Y154_SLICE_X22Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X22Y154_BO5),
.O6(CLBLM_L_X16Y154_SLICE_X22Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_L_X16Y154_SLICE_X22Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X22Y154_AO5),
.O6(CLBLM_L_X16Y154_SLICE_X22Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X23Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X23Y154_DO5),
.O6(CLBLM_L_X16Y154_SLICE_X23Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X23Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X23Y154_CO5),
.O6(CLBLM_L_X16Y154_SLICE_X23Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X23Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X23Y154_BO5),
.O6(CLBLM_L_X16Y154_SLICE_X23Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y154_SLICE_X23Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y154_SLICE_X23Y154_AO5),
.O6(CLBLM_L_X16Y154_SLICE_X23Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y125_SLICE_X2Y125_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y103_IOB_X0Y104_I),
.Q(CLBLM_R_X3Y125_SLICE_X2Y125_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafafafafafa)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y105_IOB_X0Y105_I),
.Q(CLBLM_R_X3Y126_SLICE_X2Y126_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y126_SLICE_X2Y126_AO6),
.Q(CLBLM_R_X3Y126_SLICE_X2Y126_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y126_SLICE_X2Y126_BO6),
.Q(CLBLM_R_X3Y126_SLICE_X2Y126_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303030303030)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555500000000)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_A5Q),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_F7AMUX_O),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_DO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a0a2a0a2aaa2aaa)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_CQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I3(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y131_SLICE_X1Y131_AQ),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040000044000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_BLUT (
.I0(CLBLL_L_X2Y131_SLICE_X0Y131_AO6),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I2(CLBLM_R_X3Y131_SLICE_X2Y131_CQ),
.I3(CLBLL_L_X2Y131_SLICE_X1Y131_AQ),
.I4(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I5(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf4fffff8f0fffff)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_ALUT (
.I0(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_CQ),
.I4(CLBLL_L_X2Y131_SLICE_X0Y131_BO6),
.I5(CLBLL_L_X2Y131_SLICE_X1Y131_AQ),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_BO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0022002022222020)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_DLUT (
.I0(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_DO6),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.I5(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011001011111010)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_CLUT (
.I0(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_DO6),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.I5(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3ffffffe2eeeeee)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_BLUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_DO6),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc30f3cf0d0501c50)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_ALUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_DO6),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y133_SLICE_X2Y133_AO6),
.Q(CLBLM_R_X3Y133_SLICE_X2Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777777777777)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_CLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I1(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc4cc444dddddddd)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_BLUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I2(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I3(CLBLL_L_X2Y133_SLICE_X1Y133_AQ),
.I4(CLBLL_L_X2Y132_SLICE_X1Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f3efa0f0f3efa)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_ALUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_DO6),
.I1(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I2(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c5c505f5c5c5050)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_DLUT (
.I0(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_A5Q),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555515155555551)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_CLUT (
.I0(CLBLM_R_X3Y133_SLICE_X2Y133_BO6),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_AO6),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_CO6),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200f2f022002200)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_BLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I1(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaf0aae2)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_ALUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_DO6),
.I1(CLBLL_L_X2Y131_SLICE_X0Y131_CO6),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_AO6),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_SING_X0Y199_IOB_X0Y199_I),
.Q(CLBLM_R_X3Y134_SLICE_X2Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_DO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_CO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_BO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050dc50ffffffff)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_ALUT (
.I0(LIOB33_SING_X0Y199_IOB_X0Y199_I),
.I1(CLBLL_L_X2Y131_SLICE_X0Y131_CO6),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_CO6),
.I4(CLBLL_L_X2Y131_SLICE_X0Y131_BO6),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_AO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y133_SLICE_X2Y133_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_AO5),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y133_SLICE_X2Y133_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_AO6),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y133_SLICE_X2Y133_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_BO6),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y133_SLICE_X2Y133_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_CO6),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333031)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_DLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I1(CLBLM_R_X3Y133_SLICE_X2Y133_BO5),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_DO6),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_DO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h880088008800d850)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_CLUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_CO6),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_BO5),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_CO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000500cccc0500)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_CO6),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_DO6),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.I5(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_BO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff002303aa00)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_ALUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_DO6),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_CO6),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_DO6),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_AO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y137_SLICE_X0Y137_BO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_AO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_DO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_CO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_BO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0c0c0c0c)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_AO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_DO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_CO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_BO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_AO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y137_SLICE_X2Y137_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y137_SLICE_X2Y137_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_A5Q),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y137_SLICE_X2Y137_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_CQ),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y137_SLICE_X2Y137_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafa)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_ALUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_A5Q),
.I1(1'b1),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_CQ),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_AO6),
.Q(CLBLM_R_X3Y138_SLICE_X2Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcdcdcfcfc)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_ALUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(CLBLM_R_X3Y137_SLICE_X2Y137_AO6),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y140_SLICE_X2Y140_AO5),
.Q(CLBLM_R_X3Y140_SLICE_X2Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_DO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa0aaa0aaa0aaa0)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_CLUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_CO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee000000f000f0)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_BLUT (
.I0(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I1(CLBLL_L_X2Y140_SLICE_X1Y140_AQ),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_BO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fcfc0000d278)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_ALUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_AO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_A_XOR),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_B_XOR),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_C_XOR),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_D_XOR),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y140_SLICE_X3Y140_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X3Y140_SLICE_X3Y140_D_CY, CLBLM_R_X3Y140_SLICE_X3Y140_C_CY, CLBLM_R_X3Y140_SLICE_X3Y140_B_CY, CLBLM_R_X3Y140_SLICE_X3Y140_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X3Y140_SLICE_X3Y140_DO5, CLBLM_R_X3Y140_SLICE_X2Y140_BO6, CLBLM_R_X3Y140_SLICE_X2Y140_CO6, 1'b0}),
.O({CLBLM_R_X3Y140_SLICE_X3Y140_D_XOR, CLBLM_R_X3Y140_SLICE_X3Y140_C_XOR, CLBLM_R_X3Y140_SLICE_X3Y140_B_XOR, CLBLM_R_X3Y140_SLICE_X3Y140_A_XOR}),
.S({CLBLM_R_X3Y140_SLICE_X3Y140_DO6, CLBLM_R_X3Y140_SLICE_X3Y140_CO6, CLBLM_R_X3Y140_SLICE_X3Y140_BO6, CLBLM_R_X3Y140_SLICE_X3Y140_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha9a9a5a5a5a5a5a5)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_DLUT (
.I0(CLBLL_L_X2Y140_SLICE_X1Y140_CQ),
.I1(CLBLL_L_X2Y140_SLICE_X1Y140_BQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I3(1'b1),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_DO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h669933cc6a953fc0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_CLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AO6),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I3(CLBLL_L_X2Y140_SLICE_X1Y140_BQ),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I5(CLBLL_L_X2Y140_SLICE_X1Y140_AQ),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_CO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30cfcf30659acf30)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_BLUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_AO6),
.I3(CLBLL_L_X2Y140_SLICE_X1Y140_AQ),
.I4(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_BO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_ALUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_BO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_AO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.Q(CLBLM_R_X3Y141_SLICE_X2Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaf0aaffaa00aa0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_DLUT (
.I0(CLBLM_R_X13Y147_SLICE_X19Y147_BO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ccaaccaa)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I4(CLBLM_R_X3Y141_SLICE_X2Y141_DO6),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccdcfccccc8c0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_BLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I1(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_CO6),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f500f550505050)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_DO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y141_SLICE_X3Y141_A_XOR),
.Q(CLBLM_R_X3Y141_SLICE_X3Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y141_SLICE_X3Y141_B_XOR),
.Q(CLBLM_R_X3Y141_SLICE_X3Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y141_SLICE_X3Y141_C_XOR),
.Q(CLBLM_R_X3Y141_SLICE_X3Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y141_SLICE_X3Y141_D_XOR),
.Q(CLBLM_R_X3Y141_SLICE_X3Y141_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y141_SLICE_X3Y141_CARRY4 (
.CI(CLBLM_R_X3Y140_SLICE_X3Y140_COUT),
.CO({CLBLM_R_X3Y141_SLICE_X3Y141_D_CY, CLBLM_R_X3Y141_SLICE_X3Y141_C_CY, CLBLM_R_X3Y141_SLICE_X3Y141_B_CY, CLBLM_R_X3Y141_SLICE_X3Y141_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X2Y141_SLICE_X1Y141_BQ, CLBLL_L_X2Y141_SLICE_X1Y141_AQ, CLBLL_L_X2Y140_SLICE_X1Y140_DQ, CLBLM_R_X3Y141_SLICE_X3Y141_AO5}),
.O({CLBLM_R_X3Y141_SLICE_X3Y141_D_XOR, CLBLM_R_X3Y141_SLICE_X3Y141_C_XOR, CLBLM_R_X3Y141_SLICE_X3Y141_B_XOR, CLBLM_R_X3Y141_SLICE_X3Y141_A_XOR}),
.S({CLBLM_R_X3Y141_SLICE_X3Y141_DO6, CLBLM_R_X3Y141_SLICE_X3Y141_CO6, CLBLM_R_X3Y141_SLICE_X3Y141_BO6, CLBLM_R_X3Y141_SLICE_X3Y141_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999999999999)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_DLUT (
.I0(CLBLL_L_X2Y141_SLICE_X1Y141_CQ),
.I1(CLBLL_L_X2Y141_SLICE_X1Y141_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc33cc33)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y141_SLICE_X1Y141_AQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y141_SLICE_X1Y141_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000000ffff)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X2Y140_SLICE_X1Y140_DQ),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_AQ),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0505fafafafa)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I1(1'b1),
.I2(CLBLL_L_X2Y140_SLICE_X1Y140_CQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y140_SLICE_X1Y140_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_DO6),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeaffffffff)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdfff5ff)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_CLUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfda8dd885d08dd88)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_BLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_CQ),
.I4(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I5(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaa0f000f00)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_DO6),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_AO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR),
.Q(CLBLM_R_X3Y142_SLICE_X3Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR),
.Q(CLBLM_R_X3Y142_SLICE_X3Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR),
.Q(CLBLM_R_X3Y142_SLICE_X3Y142_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR),
.Q(CLBLM_R_X3Y142_SLICE_X3Y142_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y142_SLICE_X3Y142_CARRY4 (
.CI(CLBLM_R_X3Y141_SLICE_X3Y141_COUT),
.CO({CLBLM_R_X3Y142_SLICE_X3Y142_D_CY, CLBLM_R_X3Y142_SLICE_X3Y142_C_CY, CLBLM_R_X3Y142_SLICE_X3Y142_B_CY, CLBLM_R_X3Y142_SLICE_X3Y142_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X2Y142_SLICE_X1Y142_BQ, CLBLL_L_X2Y142_SLICE_X1Y142_AQ, CLBLL_L_X2Y141_SLICE_X0Y141_AQ, CLBLL_L_X2Y141_SLICE_X1Y141_CQ}),
.O({CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR, CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR, CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR, CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR}),
.S({CLBLM_R_X3Y142_SLICE_X3Y142_DO6, CLBLM_R_X3Y142_SLICE_X3Y142_CO6, CLBLM_R_X3Y142_SLICE_X3Y142_BO6, CLBLM_R_X3Y142_SLICE_X3Y142_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0ff0f00f0f)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y142_SLICE_X1Y142_BQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y143_SLICE_X1Y143_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc33cc33)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y142_SLICE_X1Y142_AQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y142_SLICE_X1Y142_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c3c3c3c3c3c3)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y142_SLICE_X1Y142_AQ),
.I2(CLBLL_L_X2Y141_SLICE_X0Y141_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00f0f0f0f)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y141_SLICE_X0Y141_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_CQ),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3a0afa0a3a0afa0a)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I3(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8ff00f0f0ff00)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_CLUT (
.I0(CLBLM_R_X3Y137_SLICE_X2Y137_DQ),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I2(CLBLM_R_X3Y158_SLICE_X2Y158_BO6),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafad85072fa5050)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_BLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_DQ),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLL_L_X2Y158_SLICE_X0Y158_BO6),
.I5(CLBLM_R_X3Y137_SLICE_X2Y137_CQ),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf5a8a075f520a0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_ALUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I2(CLBLM_R_X3Y154_SLICE_X2Y154_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLL_L_X4Y141_SLICE_X5Y141_BQ),
.I5(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_A_XOR),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_B_XOR),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_C_XOR),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_D_XOR),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y143_SLICE_X3Y143_CARRY4 (
.CI(CLBLM_R_X3Y142_SLICE_X3Y142_COUT),
.CO({CLBLM_R_X3Y143_SLICE_X3Y143_D_CY, CLBLM_R_X3Y143_SLICE_X3Y143_C_CY, CLBLM_R_X3Y143_SLICE_X3Y143_B_CY, CLBLM_R_X3Y143_SLICE_X3Y143_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, CLBLL_L_X2Y143_SLICE_X1Y143_AQ, CLBLL_L_X2Y142_SLICE_X0Y142_AQ, CLBLL_L_X2Y143_SLICE_X1Y143_DQ}),
.O({CLBLM_R_X3Y143_SLICE_X3Y143_D_XOR, CLBLM_R_X3Y143_SLICE_X3Y143_C_XOR, CLBLM_R_X3Y143_SLICE_X3Y143_B_XOR, CLBLM_R_X3Y143_SLICE_X3Y143_A_XOR}),
.S({CLBLM_R_X3Y143_SLICE_X3Y143_DO6, CLBLM_R_X3Y143_SLICE_X3Y143_CO6, CLBLM_R_X3Y143_SLICE_X3Y143_BO6, CLBLM_R_X3Y143_SLICE_X3Y143_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999999999999)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_DLUT (
.I0(CLBLL_L_X2Y143_SLICE_X1Y143_CQ),
.I1(CLBLL_L_X2Y143_SLICE_X1Y143_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc33cc33)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y143_SLICE_X1Y143_AQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y143_SLICE_X1Y143_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c3c3c3c3c3c3)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y143_SLICE_X1Y143_AQ),
.I2(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0ff0f00f0f)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y142_SLICE_X0Y142_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y143_SLICE_X1Y143_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y144_SLICE_X2Y144_AO6),
.Q(CLBLM_R_X3Y144_SLICE_X2Y144_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffeeeffff)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_CO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I4(CLBLM_R_X3Y147_SLICE_X2Y147_DO6),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_DO6),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaaaeeaaaaaaaa)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_BO6),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f880f770fff0f)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_BLUT (
.I0(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I4(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_BO6),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_AO6),
.Q(CLBLM_R_X3Y144_SLICE_X3Y144_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000022222222)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_DLUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf05acccc)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_CLUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_BLUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_DO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe5eae04f454a40)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_BO6),
.I4(CLBLM_R_X3Y147_SLICE_X2Y147_AO6),
.I5(CLBLM_R_X3Y144_SLICE_X3Y144_CO6),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_BO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010005)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_BLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_DO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.I2(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_CO6),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0f4b0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_ALUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_BO5),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccddcccccccc)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_DLUT (
.I0(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cff0c00ccffcc00)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y158_SLICE_X3Y158_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I5(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444ccccf0f0f0f0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X3Y154_SLICE_X2Y154_AO6),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0000a202)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_ALUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_BO6),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003300130033)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_AO5),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_BO6),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_CO6),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_DO6),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1f3f3f0f3f3f3)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_CLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_AO5),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_CO6),
.I2(CLBLM_L_X10Y146_SLICE_X13Y146_CO6),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_DO6),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_CO6),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000c0c000c00)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I4(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888800330033)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_AO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_CO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0cae0cae)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffbfff)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_BLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_AO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b3a0a0a0b3a0a0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_ALUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_DLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccceecceedc)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_BO5),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00004000ccffc0ff)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffe0f0aa00aa00)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X3Y157_SLICE_X2Y157_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55fffffdfeff)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080800080800000)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_CLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_BO6),
.I5(CLBLM_R_X15Y143_SLICE_X20Y143_AO5),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040001040400000)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_BLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h007f00ff00ff00ff)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_BO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001040100000c00)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_DLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000000)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_CLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_DO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000a000a0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_BLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0f0e1f0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_ALUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heee0eeeeeeeeeeee)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_DLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_AO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.I3(CLBLM_R_X3Y148_SLICE_X3Y148_CO6),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_BO6),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000033330000)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_BO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I3(CLBLM_R_X3Y148_SLICE_X3Y148_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_CO6),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b0f080c0f0f0000)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_DLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_BO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_BO6),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff1f0fffff1f3fff)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a02000028000000)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880044444444)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_ALUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010001010100)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_DLUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000440050504400)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_CLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555557545)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I4(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500510055005100)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_DLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_AO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_CO6),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf5f555577571fff)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_CLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I1(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h90119011dbd99a9b)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_BLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333fef0f5f0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_ALUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.I2(CLBLM_R_X3Y151_SLICE_X2Y151_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000005000000044)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I3(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000320010)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_CLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I3(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000111010)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_BLUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000a0c)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_ALUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003300330023)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_DLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h050145110f09cf99)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_CLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I1(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0fff1fff5)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_BLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_DO6),
.I4(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_CO6),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff008080ff002d2d)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_ALUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I1(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_B_FDPE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h005500550000f0f0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_DLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafffffffeffffff)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_CLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I5(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f30c08f3f30c0c)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_DO5),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_CO6),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4451444003000000)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_ALUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.Q(CLBLM_R_X3Y152_SLICE_X2Y152_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f030f030b)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_BO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.I4(CLBLM_R_X3Y155_SLICE_X3Y155_CO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_BO6),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0aaaaaaa0a8a)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_CLUT (
.I0(CLBLL_L_X2Y149_SLICE_X1Y149_AO6),
.I1(CLBLL_L_X4Y156_SLICE_X4Y156_CO6),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_AO5),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_BO5),
.I5(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00cc00cc00)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_BLUT (
.I0(CLBLL_L_X2Y153_SLICE_X0Y153_DQ),
.I1(CLBLL_L_X2Y153_SLICE_X0Y153_C5Q),
.I2(1'b1),
.I3(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h550f5533ff0fff00)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_ALUT (
.I0(CLBLL_L_X2Y153_SLICE_X0Y153_DQ),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_CO6),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_AQ),
.I3(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.Q(CLBLM_R_X3Y152_SLICE_X3Y152_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffaaffbb)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_BLUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeefffffeeee)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_ALUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_CO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y153_IOB_X0Y153_I),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y153_IOB_X0Y154_I),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y155_IOB_X0Y156_I),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y157_IOB_X0Y157_I),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffaa5500)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y153_SLICE_X0Y153_A5Q),
.I3(CLBLL_L_X2Y155_SLICE_X0Y155_CO6),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_BQ),
.I5(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0055aaff)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_CLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y153_SLICE_X0Y153_AQ),
.I3(CLBLM_R_X3Y155_SLICE_X2Y155_CO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_AQ),
.I5(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000fdd0fff0fdd)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_BLUT (
.I0(CLBLM_R_X3Y157_SLICE_X3Y157_CO6),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.I2(CLBLL_L_X2Y153_SLICE_X0Y153_D5Q),
.I3(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_DQ),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8bb88cfcfcccc)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_ALUT (
.I0(CLBLL_L_X2Y153_SLICE_X0Y153_C5Q),
.I1(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_CQ),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_CO6),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y155_IOB_X0Y155_I),
.Q(CLBLM_R_X3Y153_SLICE_X3Y153_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffcc00f000cc)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y157_SLICE_X3Y157_BO6),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AQ),
.I3(CLBLL_L_X2Y152_SLICE_X0Y152_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I5(CLBLL_L_X2Y153_SLICE_X0Y153_B5Q),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.Q(CLBLM_R_X3Y154_SLICE_X2Y154_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ddf588a0dda088)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_DLUT (
.I0(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I1(CLBLM_R_X3Y154_SLICE_X2Y154_AQ),
.I2(CLBLM_R_X3Y158_SLICE_X2Y158_A5Q),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I4(CLBLM_R_X3Y155_SLICE_X2Y155_CQ),
.I5(CLBLM_R_X3Y155_SLICE_X2Y155_DQ),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_DO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f7a0a2f5d5a080)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_CLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I2(CLBLM_R_X3Y158_SLICE_X2Y158_CQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I4(CLBLM_R_X3Y154_SLICE_X2Y154_DO6),
.I5(CLBLM_R_X3Y159_SLICE_X3Y159_CQ),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_CO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2ff33e2e2cc00)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_BLUT (
.I0(CLBLM_R_X3Y155_SLICE_X2Y155_CQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I2(CLBLM_R_X3Y154_SLICE_X2Y154_AQ),
.I3(CLBLM_R_X3Y155_SLICE_X2Y155_DQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y155_SLICE_X2Y155_A5Q),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_BO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0afa0cfc0)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_ALUT (
.I0(CLBLM_R_X3Y159_SLICE_X3Y159_CQ),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_A5Q),
.I2(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I3(CLBLM_R_X3Y154_SLICE_X2Y154_BO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_AO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.Q(CLBLM_R_X3Y154_SLICE_X3Y154_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_DO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_CO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000000)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_BLUT (
.I0(CLBLM_R_X3Y157_SLICE_X3Y157_CO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_BO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_CO6),
.I4(CLBLM_R_X3Y156_SLICE_X3Y156_CO6),
.I5(CLBLL_L_X2Y155_SLICE_X0Y155_CO6),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_BO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000200)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_ALUT (
.I0(CLBLM_R_X3Y157_SLICE_X3Y157_BO6),
.I1(CLBLL_L_X2Y155_SLICE_X0Y155_BO6),
.I2(CLBLM_R_X3Y155_SLICE_X3Y155_CO6),
.I3(CLBLM_R_X3Y154_SLICE_X3Y154_BO6),
.I4(CLBLM_R_X3Y155_SLICE_X2Y155_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_AO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_A5_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y158_SLICE_X2Y158_A5Q),
.Q(CLBLM_R_X3Y155_SLICE_X2Y155_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y155_SLICE_X2Y155_AO6),
.Q(CLBLM_R_X3Y155_SLICE_X2Y155_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y154_SLICE_X2Y154_AQ),
.Q(CLBLM_R_X3Y155_SLICE_X2Y155_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y159_SLICE_X3Y159_CQ),
.Q(CLBLM_R_X3Y155_SLICE_X2Y155_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y158_SLICE_X2Y158_CQ),
.Q(CLBLM_R_X3Y155_SLICE_X2Y155_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ff55aa00)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_CQ),
.I2(CLBLM_R_X3Y155_SLICE_X2Y155_DQ),
.I3(CLBLM_R_X3Y155_SLICE_X2Y155_A5Q),
.I4(CLBLM_R_X3Y155_SLICE_X2Y155_BQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_DO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0709010e060800)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_CLUT (
.I0(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.I3(CLBLM_R_X3Y154_SLICE_X2Y154_AQ),
.I4(CLBLM_R_X3Y158_SLICE_X2Y158_A5Q),
.I5(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_CO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaafccccaaa0cccc)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_BLUT (
.I0(CLBLL_L_X2Y158_SLICE_X0Y158_CQ),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_BO6),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I5(CLBLM_R_X3Y159_SLICE_X2Y159_AQ),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_BO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y153_IOB_X0Y153_I),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_AO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y159_SLICE_X3Y159_AQ),
.Q(CLBLM_R_X3Y155_SLICE_X3Y155_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y159_SLICE_X2Y159_AQ),
.Q(CLBLM_R_X3Y155_SLICE_X3Y155_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y158_SLICE_X0Y158_CQ),
.Q(CLBLM_R_X3Y155_SLICE_X3Y155_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y155_SLICE_X2Y155_AQ),
.Q(CLBLM_R_X3Y155_SLICE_X3Y155_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfedcba9876543210)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I2(CLBLM_R_X3Y155_SLICE_X3Y155_DQ),
.I3(CLBLM_R_X3Y155_SLICE_X3Y155_AQ),
.I4(CLBLM_R_X3Y155_SLICE_X3Y155_BQ),
.I5(CLBLM_R_X3Y155_SLICE_X3Y155_CQ),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_DO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f791e680)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_CLUT (
.I0(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.I2(CLBLM_R_X3Y155_SLICE_X2Y155_AQ),
.I3(CLBLM_R_X3Y159_SLICE_X3Y159_AQ),
.I4(CLBLM_R_X3Y155_SLICE_X3Y155_DO6),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_CO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_BLUT (
.I0(CLBLM_R_X3Y159_SLICE_X3Y159_AQ),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_BQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(CLBLM_R_X3Y155_SLICE_X3Y155_CQ),
.I4(CLBLM_R_X3Y155_SLICE_X2Y155_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_BO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_ALUT (
.I0(CLBLM_R_X3Y155_SLICE_X2Y155_AQ),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_BQ),
.I2(CLBLM_R_X3Y155_SLICE_X3Y155_AQ),
.I3(CLBLM_R_X3Y155_SLICE_X3Y155_CQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_AO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y155_IOB_X0Y156_I),
.Q(CLBLM_R_X3Y156_SLICE_X2Y156_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y159_IOB_X0Y159_I),
.Q(CLBLM_R_X3Y156_SLICE_X2Y156_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y159_SLICE_X2Y159_CQ),
.Q(CLBLM_R_X3Y156_SLICE_X2Y156_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5dda0a0a088)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_DLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_BQ),
.I2(CLBLM_R_X3Y158_SLICE_X2Y158_DQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y157_SLICE_X2Y157_BO6),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_DO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccf0aa00ccf0aa)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_CLUT (
.I0(CLBLM_R_X3Y156_SLICE_X3Y156_AQ),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_CQ),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_BQ),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_CO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafbfaf8fa0b0a080)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_BLUT (
.I0(CLBLM_R_X3Y159_SLICE_X2Y159_CQ),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I2(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLM_R_X3Y158_SLICE_X2Y158_AQ),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_CO6),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_BO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f300000f0f0000)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y158_SLICE_X2Y158_AQ),
.Q(CLBLM_R_X3Y156_SLICE_X3Y156_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y155_SLICE_X1Y155_AQ),
.Q(CLBLM_R_X3Y156_SLICE_X3Y156_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y156_SLICE_X2Y156_BQ),
.Q(CLBLM_R_X3Y156_SLICE_X3Y156_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fafa5050)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_DLUT (
.I0(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I1(CLBLM_R_X3Y156_SLICE_X3Y156_CQ),
.I2(CLBLM_R_X3Y156_SLICE_X3Y156_BQ),
.I3(CLBLM_R_X3Y156_SLICE_X2Y156_CQ),
.I4(CLBLM_R_X3Y156_SLICE_X3Y156_AQ),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_DO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400041115441555)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_CLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_AQ),
.I3(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I4(CLBLM_R_X3Y156_SLICE_X3Y156_DO6),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_BQ),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_CO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffaaf0cc00aaf0)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_BLUT (
.I0(CLBLM_R_X3Y156_SLICE_X3Y156_AQ),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_AQ),
.I2(CLBLM_R_X3Y156_SLICE_X3Y156_CQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_CQ),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_BO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5702fda85500)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_ALUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(CLBLM_R_X3Y156_SLICE_X3Y156_BO6),
.I4(CLBLM_R_X3Y158_SLICE_X2Y158_AQ),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_BQ),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y155_IOB_X0Y155_I),
.Q(CLBLM_R_X3Y157_SLICE_X2Y157_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y157_IOB_X0Y157_I),
.Q(CLBLM_R_X3Y157_SLICE_X2Y157_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y158_SLICE_X2Y158_BQ),
.Q(CLBLM_R_X3Y157_SLICE_X2Y157_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y158_SLICE_X2Y158_DQ),
.Q(CLBLM_R_X3Y157_SLICE_X2Y157_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_DO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_CO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_BLUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_BQ),
.I1(CLBLM_R_X3Y157_SLICE_X2Y157_DQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(CLBLM_R_X3Y157_SLICE_X2Y157_CQ),
.I4(CLBLM_R_X3Y157_SLICE_X3Y157_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_BO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88fc3000000000)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_ALUT (
.I0(CLBLM_R_X3Y157_SLICE_X3Y157_AQ),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I2(CLBLM_R_X3Y157_SLICE_X3Y157_AO6),
.I3(CLBLM_R_X3Y158_SLICE_X2Y158_BQ),
.I4(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_BO6),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y165_IOB_X0Y165_I),
.Q(CLBLM_R_X3Y157_SLICE_X3Y157_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y171_IOB_X0Y172_I),
.Q(CLBLM_R_X3Y157_SLICE_X3Y157_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y157_SLICE_X3Y157_AQ),
.Q(CLBLM_R_X3Y157_SLICE_X3Y157_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y157_SLICE_X2Y157_BQ),
.Q(CLBLM_R_X3Y157_SLICE_X3Y157_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccaaf000ccaaf0)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_DLUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_CQ),
.I1(CLBLM_R_X3Y157_SLICE_X3Y157_CQ),
.I2(CLBLM_R_X3Y157_SLICE_X3Y157_DQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y157_SLICE_X2Y157_DQ),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_DO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddf888addd58880)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_CLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I1(CLBLM_R_X3Y157_SLICE_X3Y157_AQ),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I4(CLBLM_R_X3Y157_SLICE_X3Y157_DO6),
.I5(CLBLM_R_X3Y157_SLICE_X2Y157_BQ),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_CO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0c03000e020e02)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_BLUT (
.I0(CLBLM_R_X3Y158_SLICE_X3Y158_DO6),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.I3(CLBLM_R_X3Y159_SLICE_X3Y159_BQ),
.I4(CLBLM_R_X3Y157_SLICE_X2Y157_AQ),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_BO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33b8b8cc00b8b8)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_ALUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_DQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I2(CLBLM_R_X3Y157_SLICE_X3Y157_CQ),
.I3(CLBLM_R_X3Y157_SLICE_X2Y157_BQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y157_SLICE_X2Y157_CQ),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_AO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_A5_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y157_IOB_X0Y158_I),
.Q(CLBLM_R_X3Y158_SLICE_X2Y158_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y158_SLICE_X2Y158_AO6),
.Q(CLBLM_R_X3Y158_SLICE_X2Y158_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y173_IOB_X0Y173_I),
.Q(CLBLM_R_X3Y158_SLICE_X2Y158_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y173_IOB_X0Y174_I),
.Q(CLBLM_R_X3Y158_SLICE_X2Y158_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y181_IOB_X0Y181_I),
.Q(CLBLM_R_X3Y158_SLICE_X2Y158_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_DO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_CO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0dd88f0f0)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLM_R_X3Y159_SLICE_X2Y159_DQ),
.I2(CLBLM_R_X3Y158_SLICE_X3Y158_CO6),
.I3(CLBLM_R_X3Y159_SLICE_X2Y159_BQ),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_BO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y167_IOB_X0Y167_I),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y159_SLICE_X3Y159_BQ),
.Q(CLBLM_R_X3Y158_SLICE_X3Y158_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y159_SLICE_X2Y159_BQ),
.Q(CLBLM_R_X3Y158_SLICE_X3Y158_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y159_SLICE_X2Y159_DQ),
.Q(CLBLM_R_X3Y158_SLICE_X3Y158_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y157_SLICE_X2Y157_AQ),
.Q(CLBLM_R_X3Y158_SLICE_X3Y158_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888fc30fc30)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_DLUT (
.I0(CLBLM_R_X3Y158_SLICE_X3Y158_CQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I2(CLBLM_R_X3Y158_SLICE_X3Y158_DQ),
.I3(CLBLM_R_X3Y158_SLICE_X3Y158_BQ),
.I4(CLBLM_R_X3Y158_SLICE_X3Y158_AQ),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_DO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaccccf0f0)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_CLUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_AQ),
.I1(CLBLM_R_X3Y158_SLICE_X3Y158_CQ),
.I2(CLBLM_R_X3Y158_SLICE_X3Y158_BQ),
.I3(CLBLM_R_X3Y159_SLICE_X3Y159_BQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_CO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd855d8aad800d8)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLM_R_X3Y158_SLICE_X3Y158_BQ),
.I2(CLBLM_R_X3Y158_SLICE_X3Y158_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I4(CLBLM_R_X3Y157_SLICE_X2Y157_AQ),
.I5(CLBLM_R_X3Y158_SLICE_X3Y158_CQ),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_BO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff1ff010ef0fe000)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_AQ),
.I2(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I3(CLBLM_R_X3Y159_SLICE_X2Y159_BQ),
.I4(CLBLM_R_X3Y158_SLICE_X3Y158_BO6),
.I5(CLBLM_R_X3Y159_SLICE_X3Y159_BQ),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_AO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y159_SLICE_X2Y159_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y169_IOB_X0Y169_I),
.Q(CLBLM_R_X3Y159_SLICE_X2Y159_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y159_SLICE_X2Y159_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y171_IOB_X0Y171_I),
.Q(CLBLM_R_X3Y159_SLICE_X2Y159_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y159_SLICE_X2Y159_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y175_IOB_X0Y175_I),
.Q(CLBLM_R_X3Y159_SLICE_X2Y159_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y159_SLICE_X2Y159_D_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y179_IOB_X0Y179_I),
.Q(CLBLM_R_X3Y159_SLICE_X2Y159_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y159_SLICE_X2Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y159_SLICE_X2Y159_DO5),
.O6(CLBLM_R_X3Y159_SLICE_X2Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y159_SLICE_X2Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y159_SLICE_X2Y159_CO5),
.O6(CLBLM_R_X3Y159_SLICE_X2Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y159_SLICE_X2Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y159_SLICE_X2Y159_BO5),
.O6(CLBLM_R_X3Y159_SLICE_X2Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y159_SLICE_X2Y159_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y159_SLICE_X2Y159_AO5),
.O6(CLBLM_R_X3Y159_SLICE_X2Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y159_SLICE_X3Y159_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y161_IOB_X0Y161_I),
.Q(CLBLM_R_X3Y159_SLICE_X3Y159_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y159_SLICE_X3Y159_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y163_IOB_X0Y163_I),
.Q(CLBLM_R_X3Y159_SLICE_X3Y159_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y159_SLICE_X3Y159_C_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_X0Y165_IOB_X0Y166_I),
.Q(CLBLM_R_X3Y159_SLICE_X3Y159_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y159_SLICE_X3Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y159_SLICE_X3Y159_DO5),
.O6(CLBLM_R_X3Y159_SLICE_X3Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y159_SLICE_X3Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y159_SLICE_X3Y159_CO5),
.O6(CLBLM_R_X3Y159_SLICE_X3Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y159_SLICE_X3Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y159_SLICE_X3Y159_BO5),
.O6(CLBLM_R_X3Y159_SLICE_X3Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y159_SLICE_X3Y159_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y159_SLICE_X3Y159_AO5),
.O6(CLBLM_R_X3Y159_SLICE_X3Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0503050305030503)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0afcfaccaaccaa)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_BLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0e4ffcc00cc)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_ALUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y128_SLICE_X7Y128_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X5Y128_SLICE_X7Y128_D_CY, CLBLM_R_X5Y128_SLICE_X7Y128_C_CY, CLBLM_R_X5Y128_SLICE_X7Y128_B_CY, CLBLM_R_X5Y128_SLICE_X7Y128_A_CY}),
.CYINIT(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.DI({1'b0, 1'b0, 1'b0, CLBLM_R_X5Y128_SLICE_X7Y128_AO5}),
.O({CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR, CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR, CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR, CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR}),
.S({CLBLM_R_X5Y128_SLICE_X7Y128_DO6, CLBLM_R_X5Y128_SLICE_X7Y128_CO6, CLBLM_R_X5Y128_SLICE_X7Y128_BO6, CLBLM_R_X5Y128_SLICE_X7Y128_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_BO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_CO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_DO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55cfcfcf55c0c0c0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_DLUT (
.I0(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55fc550cfcfc0c0c)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_CLUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h54fe04aefcfc0c0c)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_BLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I3(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeba5410fc30fc30)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_ALUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y129_SLICE_X7Y129_CARRY4 (
.CI(CLBLM_R_X5Y128_SLICE_X7Y128_COUT),
.CO({CLBLM_R_X5Y129_SLICE_X7Y129_D_CY, CLBLM_R_X5Y129_SLICE_X7Y129_C_CY, CLBLM_R_X5Y129_SLICE_X7Y129_B_CY, CLBLM_R_X5Y129_SLICE_X7Y129_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR, CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR, CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR, CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR}),
.S({CLBLM_R_X5Y129_SLICE_X7Y129_DO6, CLBLM_R_X5Y129_SLICE_X7Y129_CO6, CLBLM_R_X5Y129_SLICE_X7Y129_BO6, CLBLM_R_X5Y129_SLICE_X7Y129_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X5Y130_SLICE_X6Y130_D_CY, CLBLM_R_X5Y130_SLICE_X6Y130_C_CY, CLBLM_R_X5Y130_SLICE_X6Y130_B_CY, CLBLM_R_X5Y130_SLICE_X6Y130_A_CY}),
.CYINIT(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.DI({1'b0, 1'b0, 1'b0, CLBLM_R_X5Y130_SLICE_X6Y130_AO5}),
.O({CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR, CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR, CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR, CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR}),
.S({CLBLM_R_X5Y130_SLICE_X6Y130_DO6, CLBLM_R_X5Y130_SLICE_X6Y130_CO6, CLBLM_R_X5Y130_SLICE_X6Y130_BO6, CLBLM_R_X5Y130_SLICE_X6Y130_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CARRY4 (
.CI(CLBLM_R_X5Y129_SLICE_X7Y129_COUT),
.CO({CLBLM_R_X5Y130_SLICE_X7Y130_D_CY, CLBLM_R_X5Y130_SLICE_X7Y130_C_CY, CLBLM_R_X5Y130_SLICE_X7Y130_B_CY, CLBLM_R_X5Y130_SLICE_X7Y130_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR, CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR, CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR, CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR}),
.S({CLBLM_R_X5Y130_SLICE_X7Y130_DO6, CLBLM_R_X5Y130_SLICE_X7Y130_CO6, CLBLM_R_X5Y130_SLICE_X7Y130_BO6, CLBLM_R_X5Y130_SLICE_X7Y130_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y131_SLICE_X6Y131_CARRY4 (
.CI(CLBLM_R_X5Y130_SLICE_X6Y130_COUT),
.CO({CLBLM_R_X5Y131_SLICE_X6Y131_D_CY, CLBLM_R_X5Y131_SLICE_X6Y131_C_CY, CLBLM_R_X5Y131_SLICE_X6Y131_B_CY, CLBLM_R_X5Y131_SLICE_X6Y131_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR, CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR, CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR, CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR}),
.S({CLBLM_R_X5Y131_SLICE_X6Y131_DO6, CLBLM_R_X5Y131_SLICE_X6Y131_CO6, CLBLM_R_X5Y131_SLICE_X6Y131_BO6, CLBLM_R_X5Y131_SLICE_X6Y131_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y131_SLICE_X7Y131_CARRY4 (
.CI(CLBLM_R_X5Y130_SLICE_X7Y130_COUT),
.CO({CLBLM_R_X5Y131_SLICE_X7Y131_D_CY, CLBLM_R_X5Y131_SLICE_X7Y131_C_CY, CLBLM_R_X5Y131_SLICE_X7Y131_B_CY, CLBLM_R_X5Y131_SLICE_X7Y131_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y131_SLICE_X7Y131_D_XOR, CLBLM_R_X5Y131_SLICE_X7Y131_C_XOR, CLBLM_R_X5Y131_SLICE_X7Y131_B_XOR, CLBLM_R_X5Y131_SLICE_X7Y131_A_XOR}),
.S({CLBLM_R_X5Y131_SLICE_X7Y131_DO6, CLBLM_R_X5Y131_SLICE_X7Y131_CO6, CLBLM_R_X5Y131_SLICE_X7Y131_BO6, CLBLM_R_X5Y131_SLICE_X7Y131_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y132_SLICE_X6Y132_CARRY4 (
.CI(CLBLM_R_X5Y131_SLICE_X6Y131_COUT),
.CO({CLBLM_R_X5Y132_SLICE_X6Y132_D_CY, CLBLM_R_X5Y132_SLICE_X6Y132_C_CY, CLBLM_R_X5Y132_SLICE_X6Y132_B_CY, CLBLM_R_X5Y132_SLICE_X6Y132_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR, CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR, CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR, CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR}),
.S({CLBLM_R_X5Y132_SLICE_X6Y132_DO6, CLBLM_R_X5Y132_SLICE_X6Y132_CO6, CLBLM_R_X5Y132_SLICE_X6Y132_BO6, CLBLM_R_X5Y132_SLICE_X6Y132_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h001d001dff1dff1d)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_A_CY),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_D_CY),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8fcfc3030fcfc30)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_CO6),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h44eeeeee44ee4444)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_CO6),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I2(1'b1),
.I3(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00001155000030f0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_ALUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I5(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y133_SLICE_X6Y133_CARRY4 (
.CI(CLBLM_R_X5Y132_SLICE_X6Y132_COUT),
.CO({CLBLM_R_X5Y133_SLICE_X6Y133_D_CY, CLBLM_R_X5Y133_SLICE_X6Y133_C_CY, CLBLM_R_X5Y133_SLICE_X6Y133_B_CY, CLBLM_R_X5Y133_SLICE_X6Y133_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y133_SLICE_X6Y133_D_XOR, CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR, CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR, CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR}),
.S({CLBLM_R_X5Y133_SLICE_X6Y133_DO6, CLBLM_R_X5Y133_SLICE_X6Y133_CO6, CLBLM_R_X5Y133_SLICE_X6Y133_BO6, CLBLM_R_X5Y133_SLICE_X6Y133_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_BO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_DLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I4(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I5(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f005f508f80dfd)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.I3(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_BO6),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ccffcc00acffac)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_BO6),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7373ff7351515151)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I3(CLBLL_L_X2Y131_SLICE_X0Y131_CO6),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_CO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaee222a2aee22)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_DO6),
.I3(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccee4ecccc444e)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_BLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.I2(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_CO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fa50f0f07272)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_ALUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X8Y138_SLICE_X11Y138_BO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaea2aea2)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_DLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_BO6),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fdff2000)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffdd88008800)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_BLUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefc00001030)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_ALUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_DO6),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_AO6),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_CO6),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_BO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a00020000000000)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fffdfff0fffcfff)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_CLUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h45ef44ee40ea44ee)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_BLUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.I3(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050fbea5140)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_ALUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_CO6),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000ffff)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.I5(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33fff3ffbbfffbff)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22220000ffff5555)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I1(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000d8fff0ffd8)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I3(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_AO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_BO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f7fff7f7f7fff7)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_CO6),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7f7700000000)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_DO6),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0cceef0f0cc44)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f0e4f0a0f0e4)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_DO6),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_BO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_CO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_D_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_DO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f088f0ddf0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_DLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_DQ),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_CO6),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0cccccfc5cccc)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I5(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffd2220dfdd0200)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_BLUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_DO6),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X13Y147_SLICE_X19Y147_BO6),
.I4(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000fff1d111ddd)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_ALUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I2(LIOB33_X0Y189_IOB_X0Y189_I),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I4(CLBLM_R_X5Y136_SLICE_X7Y136_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_DO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7ffffff777ffff)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_AO5),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_BO6),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fdfffff5fdf5f5f)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_CLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_BO6),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heee4eecc44e444cc)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_CO6),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f00df800000cccc)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_ALUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_BO6),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_CO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000e2e20000f3c0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_DLUT (
.I0(CLBLM_R_X15Y140_SLICE_X21Y140_DO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffb00c8ff730040)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_CO6),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f55550f335533)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_BLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I2(LIOB33_X0Y181_IOB_X0Y182_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f55550f335533)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I2(LIOB33_X0Y183_IOB_X0Y184_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1515151505550050)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_DLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_AO6),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I3(CLBLM_R_X15Y143_SLICE_X21Y143_AO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb8bbbbb88b88888)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_CO6),
.I4(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I5(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fffff3f1)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_BLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_BO6),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_AO6),
.I3(CLBLM_R_X15Y143_SLICE_X21Y143_AO6),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_AO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_AO5),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f0f4f0f050f050)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_CO5),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5a0a0a0a0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I1(1'b1),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11f0f0bb11bb11)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_CLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I1(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.I3(CLBLM_R_X7Y138_SLICE_X8Y138_C_XOR),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccceeee00cc0000)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_BLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0300000aa33aa33)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_ALUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_B_XOR),
.I1(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_AO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffdfffffffffff)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_DLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_CO6),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500ffaadf80)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5000000f7333333)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_BLUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_CQ),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_BO6),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_R_X5Y139_SLICE_X6Y139_CO6),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X13Y141_SLICE_X19Y141_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO5),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff7fffff)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_CLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_CO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb070000080400000)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_BLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_DO6),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff2000005555ffff)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5ffffffffffff)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff5ffff7777ffff)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_DO6),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf870f870f0f0f0f0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_ALUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_AO5),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_BO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_CO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f099f0aa)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_DLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_CO6),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.I4(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hea2aaaaaea2aaaaa)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_CLUT (
.I0(CLBLM_R_X13Y147_SLICE_X19Y147_BO6),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44cccccccccccc)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_BLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_BO6),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66006600f8f070f0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_ALUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I2(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_CO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacff00acacff00)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_BLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_DO6),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7e69180f7e69180)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_DO6),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_AO6),
.I4(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X5Y141_SLICE_X6Y141_MUXF7A (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_BO6),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_AO6),
.O(CLBLM_R_X5Y141_SLICE_X6Y141_F7AMUX_O),
.S(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_CO6),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5aff006666ff00)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_DLUT (
.I0(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaa0aaaaaaaaaaa)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_CLUT (
.I0(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacfcfcacac0c0c)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_BLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_BO6),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdf8585dada8080)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.I5(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X5Y141_SLICE_X7Y141_MUXF7A (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_BO6),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.O(CLBLM_R_X5Y141_SLICE_X7Y141_F7AMUX_O),
.S(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y142_SLICE_X6Y142_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X5Y142_SLICE_X6Y142_D_CY, CLBLM_R_X5Y142_SLICE_X6Y142_C_CY, CLBLM_R_X5Y142_SLICE_X6Y142_B_CY, CLBLM_R_X5Y142_SLICE_X6Y142_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X3Y140_SLICE_X3Y140_DQ, CLBLM_R_X3Y140_SLICE_X3Y140_CQ, CLBLM_R_X3Y140_SLICE_X3Y140_BQ, CLBLM_R_X3Y140_SLICE_X3Y140_AQ}),
.O({CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR, CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR, CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR, CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR}),
.S({CLBLM_R_X5Y142_SLICE_X6Y142_DO6, CLBLM_R_X5Y142_SLICE_X6Y142_CO6, CLBLM_R_X5Y142_SLICE_X6Y142_BO6, CLBLM_R_X5Y142_SLICE_X6Y142_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9933993399cc99cc)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_DLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_BO6),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0af55fa00af55fa0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ccc3c333ccc3c3)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.I3(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c0f3c0f3cf03cf0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cafa0afa0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_DLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bb88bb88)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222ee22ee22)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_DO6),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55bbbbaa001111)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I5(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X5Y142_SLICE_X7Y142_MUXF7A (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_AO6),
.O(CLBLM_R_X5Y142_SLICE_X7Y142_F7AMUX_O),
.S(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y143_SLICE_X6Y143_CARRY4 (
.CI(CLBLM_R_X5Y142_SLICE_X6Y142_COUT),
.CO({CLBLM_R_X5Y143_SLICE_X6Y143_D_CY, CLBLM_R_X5Y143_SLICE_X6Y143_C_CY, CLBLM_R_X5Y143_SLICE_X6Y143_B_CY, CLBLM_R_X5Y143_SLICE_X6Y143_A_CY}),
.CYINIT(1'b0),
.DI({CLBLM_R_X3Y141_SLICE_X3Y141_DQ, CLBLM_R_X3Y141_SLICE_X3Y141_CQ, CLBLM_R_X3Y141_SLICE_X3Y141_BQ, CLBLM_R_X3Y141_SLICE_X3Y141_AQ}),
.O({CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR, CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR, CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR, CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR}),
.S({CLBLM_R_X5Y143_SLICE_X6Y143_DO6, CLBLM_R_X5Y143_SLICE_X6Y143_CO6, CLBLM_R_X5Y143_SLICE_X6Y143_BO6, CLBLM_R_X5Y143_SLICE_X6Y143_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y141_SLICE_X3Y141_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf50af5005fa05fa)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_DO6),
.I3(CLBLM_R_X3Y141_SLICE_X3Y141_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cc3333cccccc)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y141_SLICE_X3Y141_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_CO6),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f3c0f3cf03cf03c)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_BO6),
.I2(CLBLM_R_X3Y141_SLICE_X3Y141_AQ),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ee44ee44ee44ee4)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.I3(CLBLM_R_X5Y145_SLICE_X7Y145_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcccccecececec)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_CLUT (
.I0(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.I1(CLBLL_L_X4Y145_SLICE_X5Y145_AO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_DO6),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3fcc0cf333c000)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_CO6),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf791e680f791e680)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X5Y143_SLICE_X7Y143_MUXF7A (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_AO6),
.O(CLBLM_R_X5Y143_SLICE_X7Y143_F7AMUX_O),
.S(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y144_SLICE_X6Y144_CARRY4 (
.CI(CLBLM_R_X5Y143_SLICE_X6Y143_COUT),
.CO({CLBLM_R_X5Y144_SLICE_X6Y144_D_CY, CLBLM_R_X5Y144_SLICE_X6Y144_C_CY, CLBLM_R_X5Y144_SLICE_X6Y144_B_CY, CLBLM_R_X5Y144_SLICE_X6Y144_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y144_SLICE_X6Y144_D_XOR, CLBLM_R_X5Y144_SLICE_X6Y144_C_XOR, CLBLM_R_X5Y144_SLICE_X6Y144_B_XOR, CLBLM_R_X5Y144_SLICE_X6Y144_A_XOR}),
.S({CLBLM_R_X5Y144_SLICE_X6Y144_DO6, CLBLM_R_X5Y144_SLICE_X6Y144_CO6, CLBLM_R_X5Y144_SLICE_X6Y144_BO6, CLBLM_R_X5Y144_SLICE_X6Y144_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7d7d7d28282828)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_AO6),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_CLUT (
.I0(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_BO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_DO6),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff1111111f111111)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_BLUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_DO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00000000101)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000003)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_ALUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_DQ),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_A_CY),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_BO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f000f000f)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeeeef0f0f0f0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I4(CLBLL_L_X4Y151_SLICE_X5Y151_AO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff3070)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_AO6),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03130303ffaa0000)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_BO6),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffcc00ccf5cc)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_CLUT (
.I0(CLBLM_R_X5Y151_SLICE_X7Y151_AO5),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_DO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_DO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500330033)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffafff88ff8c)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_ALUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_DO6),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_BO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffe0f3ffff)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_DLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040000000080)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888c8880888880)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_BO5),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0f0c0d0c)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_ALUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_DO6),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_CO6),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff1fff1ff31ff31)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_AO5),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_CO6),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_AO6),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1011101011111111)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_BLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_CO6),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I3(CLBLM_R_X7Y148_SLICE_X9Y148_BO6),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_AO6),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff7fff5fff5fff)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I3(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000800000)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_DLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_BO6),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3faaffaaffaaffaa)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X7Y148_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffee44444444)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_BLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffacccccffc)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_ALUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_CO6),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7030c0c07030f0f0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_CO6),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h110800003f080000)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f500f500f500e4)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_BLUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_DO6),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_CO6),
.I2(CLBLM_L_X16Y142_SLICE_X22Y142_AO5),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_CO6),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_AO5),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400050440415)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_AO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haabaaaaaaaaaabaa)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_DLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_BO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000888c0000800c)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I5(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefcfffffffff)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_BLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff2323ffff2223)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_DO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_DO6),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_BO6),
.I4(CLBLM_R_X5Y151_SLICE_X7Y151_CO6),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_CO6),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000000000000)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_CLUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.I5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0bfaf00003300)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202020222a22222)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_AO6),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f00aaaabdbb)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc000000c080)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa5555ffff3333)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fcfd0000fcfc)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_ALUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_DO5),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_BO6),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_AO6),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_BO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f060a0b)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_BO6),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000042420206)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_CLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe7e7ffffffaaff)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_BLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc0ccc0c)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0305020002000244)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05550000cdddcccc)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_CLUT (
.I0(CLBLM_R_X5Y151_SLICE_X7Y151_AO6),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLM_R_X5Y151_SLICE_X7Y151_DO6),
.I5(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffbffffff)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I3(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7fffcfcfcf0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_ALUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbb8b88b8b8888)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_BLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f00fff0fff0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_BO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffffffffff)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_DLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd555aaaa5555aaaa)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7df5f5f5c0000000)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f3d1f3c0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BO6),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_CO6),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa00000000)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_DLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00000000000000)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haffa000023320000)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_DO6),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacfc0cfc0cfc0cf)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_DO6),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd0ddd0ffff0000)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_BLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ff00f0f0f0f0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_ALUT (
.I0(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I1(1'b1),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_CO6),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaffaa00aa00aa)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_DLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_DQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_BO6),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he666cccc80000000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_BLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3aff3aff3a003a00)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_ALUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_DO6),
.I1(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555500000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_ALUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c3f11110c3fdddd)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff04f700ff15d5)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_BLUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333313b3237303f)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1105bb0511afbbaf)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_BLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333312033333b7f)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505f5f03f303f3)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c3f3f11dd11dd)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_DQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_CQ),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h330f0055330fff55)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_BLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a044004400)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555505000000000)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_AQ),
.I3(1'b1),
.I4(CLBLM_L_X16Y136_SLICE_X22Y136_BQ),
.I5(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555553535533)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_CLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100fdff0111fddd)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_BLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h01555555fc000000)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_DO6),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_AQ),
.I2(CLBLM_L_X16Y136_SLICE_X22Y136_BQ),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111dddddd11dd11)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_DLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I2(1'b1),
.I3(CLBLL_L_X26Y136_SLICE_X38Y136_AO5),
.I4(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3301332300010023)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_CLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_AO5),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I4(CLBLM_R_X7Y135_SLICE_X8Y135_DO6),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h051105bbaf11afbb)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.I2(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaafaf00004400)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_AO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_BO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h75ffffff30ffffff)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_DLUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0000000880088)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I1(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_DO6),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_BO6),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555cfc05555cccc)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_BLUT (
.I0(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555f0f05555ccf0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_ALUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I3(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55335533f033f033)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0055aaff)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_CLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_BO5),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_DO6),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfef7fdbfef7fdf)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_BLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f0f0e2e2f0f0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_ALUT (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.I2(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000408000400)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_CO6),
.I2(CLBLM_R_X7Y136_SLICE_X8Y136_BO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffff7ff)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_CLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8fa88aaf8f08800)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_F8MUX_O),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_DO6),
.I5(CLBLM_R_X11Y137_SLICE_X14Y137_F8MUX_O),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ffaa00aa)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_ALUT (
.I0(CLBLM_R_X7Y137_SLICE_X9Y137_DO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_CO6),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303f3fafa0afa0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_DLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_AO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffd0020fff80070)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_AO6),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_BO6),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe5ef454ae0ea404)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_BLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_AQ),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I5(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7e6b3a2d5c49180)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_ALUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.I3(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X7Y137_SLICE_X8Y137_MUXF7A (
.I0(CLBLM_R_X7Y137_SLICE_X8Y137_BO6),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.O(CLBLM_R_X7Y137_SLICE_X8Y137_F7AMUX_O),
.S(CLBLM_R_X5Y137_SLICE_X7Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc307777fc304444)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_AO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I3(CLBLM_L_X16Y137_SLICE_X22Y137_BO5),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d855ffd8d800aa)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I1(CLBLM_R_X13Y137_SLICE_X19Y137_AO5),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I5(CLBLL_L_X4Y137_SLICE_X5Y137_AQ),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1f0e0f0fbf040)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_BLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_AO6),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h53ff530f0000ffff)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.I1(CLBLM_R_X15Y140_SLICE_X21Y140_AO5),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X7Y138_SLICE_X8Y138_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X7Y138_SLICE_X8Y138_D_CY, CLBLM_R_X7Y138_SLICE_X8Y138_C_CY, CLBLM_R_X7Y138_SLICE_X8Y138_B_CY, CLBLM_R_X7Y138_SLICE_X8Y138_A_CY}),
.CYINIT(CLBLM_R_X5Y138_SLICE_X7Y138_DO6),
.DI({CLBLM_R_X5Y140_SLICE_X6Y140_CO6, CLBLM_R_X5Y140_SLICE_X6Y140_CO6, CLBLM_R_X5Y140_SLICE_X6Y140_CO6, CLBLM_R_X7Y138_SLICE_X8Y138_AO5}),
.O({CLBLM_R_X7Y138_SLICE_X8Y138_D_XOR, CLBLM_R_X7Y138_SLICE_X8Y138_C_XOR, CLBLM_R_X7Y138_SLICE_X8Y138_B_XOR, CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR}),
.S({CLBLM_R_X7Y138_SLICE_X8Y138_DO6, CLBLM_R_X7Y138_SLICE_X8Y138_CO6, CLBLM_R_X7Y138_SLICE_X8Y138_BO6, CLBLM_R_X7Y138_SLICE_X8Y138_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555333355a533c3)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_DLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I1(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010ef10efefef10)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_CLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I3(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I5(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300ffcc390af5c6)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I3(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f8f0f0ff77ffff)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_AO5),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30000300c0000c00)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_CO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0104020810402080)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_CLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0015551500105510)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_BLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I1(CLBLM_R_X13Y141_SLICE_X19Y141_CO6),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_AO6),
.I5(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h725072faccffcc00)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_D_XOR),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X7Y139_SLICE_X8Y139_CARRY4 (
.CI(CLBLM_R_X7Y138_SLICE_X8Y138_COUT),
.CO({CLBLM_R_X7Y139_SLICE_X8Y139_D_CY, CLBLM_R_X7Y139_SLICE_X8Y139_C_CY, CLBLM_R_X7Y139_SLICE_X8Y139_B_CY, CLBLM_R_X7Y139_SLICE_X8Y139_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, CLBLM_R_X5Y140_SLICE_X6Y140_CO6, CLBLM_R_X5Y140_SLICE_X6Y140_CO6, CLBLM_R_X5Y140_SLICE_X6Y140_CO6}),
.O({CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR, CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR, CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR, CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR}),
.S({CLBLM_R_X7Y139_SLICE_X8Y139_DO6, CLBLM_R_X7Y139_SLICE_X8Y139_CO6, CLBLM_R_X7Y139_SLICE_X8Y139_BO6, CLBLM_R_X7Y139_SLICE_X8Y139_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h74747474748b7474)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_DLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50635050fac9fafa)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_CLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333f0f03399f05a)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_CQ),
.I2(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffcccc0af5c6c6)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h555500ff0f0f0f0f)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_DLUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR),
.I1(1'b1),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I3(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03034477cfcf4477)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_CLUT (
.I0(CLBLM_R_X15Y142_SLICE_X20Y142_BO6),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000c5c5c5c5)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_BLUT (
.I0(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I3(CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5cccca0f5a0f5)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_ALUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.I2(CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000880000f0f8)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_DO6),
.I2(CLBLM_R_X11Y137_SLICE_X15Y137_AO5),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_F7AMUX_O),
.I5(CLBLM_R_X7Y140_SLICE_X8Y140_BO6),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffffffffffff)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_BLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff20ff00ffffff00)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_BO6),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_DO6),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_DO6),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_CO6),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_CO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005000000050505)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_DLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_F7AMUX_O),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_F7AMUX_O),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333303000302)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_CLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_AO6),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_CO6),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_BO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.I5(CLBLM_R_X7Y140_SLICE_X8Y140_AO6),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cafafa0a0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_BLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe3ece0ef232c202)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X7Y140_SLICE_X9Y140_MUXF7A (
.I0(CLBLM_R_X7Y140_SLICE_X9Y140_BO6),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_AO6),
.O(CLBLM_R_X7Y140_SLICE_X9Y140_F7AMUX_O),
.S(CLBLM_R_X5Y137_SLICE_X7Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3344cc3f3377cc3f)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_DLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_AO5),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffddfffffffdff)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd111130fc30fc)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_BLUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I3(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d001d331dcc1dff)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_ALUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I4(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I5(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X7Y141_SLICE_X8Y141_MUXF7A (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_BO6),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_AO6),
.O(CLBLM_R_X7Y141_SLICE_X8Y141_F7AMUX_O),
.S(CLBLM_R_X5Y137_SLICE_X7Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1f3e2c0f3f3c0c0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_DLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_CQ),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_CO6),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeaaabfffeaffbf)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_CLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_CQ),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_CO6),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.I5(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf5fffff3f5fffff)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_BLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_CQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_CO6),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ffbfbf00bf)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_BO6),
.I4(CLBLM_R_X5Y139_SLICE_X7Y139_AO6),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO5),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101232311331133)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLM_R_X15Y139_SLICE_X21Y139_AO5),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_AO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaf3323ffff3333)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_CO6),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_AO6),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ec00cc00cc00)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO5),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000faffffff)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_BO6),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f000b000)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_CLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_BO6),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555577775fff)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_DO6),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555547748bb8)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_BO6),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fff40004000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_BLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I4(1'b1),
.I5(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaa2aaa30003000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_ALUT (
.I0(CLBLM_R_X15Y148_SLICE_X21Y148_BO6),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I4(CLBLM_R_X11Y145_SLICE_X15Y145_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff505f00ff00ff)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_BLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c0ffff0000ffff)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbfffb)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_AO5),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heefaeefaffaa00aa)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_BQ),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f0000fffffcff)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_CO6),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff007700ff003f00)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_ALUT (
.I0(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_BO6),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I5(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ff55aa00)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_DLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I3(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_DO6),
.I5(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h082a193b4c6e5d7f)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_DO6),
.I5(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaeff00afaaff00)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_BLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff33330f0f5555)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_DO6),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacac00000055)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_BLUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_A_CY),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30eeee2222)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_ALUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddd88888888)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefe44dceedc44)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_CLUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_DQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I4(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0ffa0ff00000044)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_BLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_BO6),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I5(CLBLM_R_X7Y145_SLICE_X9Y145_CO6),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0aaf0aa)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_ALUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I4(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabaaaaaaabfeaaa)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffa0df08f7)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbeafbeafbfbaaaa)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_BO6),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_CO5),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_AO5),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc30b8fcfc30fc)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_BLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_DO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I4(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_CO6),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccefeeefef)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_DO6),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_CO6),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AO6),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff773232)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100000000000)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdfff)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0077003300550000)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_DO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I4(CLBLM_L_X8Y149_SLICE_X10Y149_CO5),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_DO6),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100330133)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_DLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_CO6),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.I4(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0dd333a040a040)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000ffffaaaa)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcccfccc0fffffff)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f2f8f0f88228800)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_DLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddfddffffffffef)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_BO5),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000222200000000)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00400004ffdffff7)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h050000a308080c00)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffff08080808)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_BLUT (
.I0(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5510555045000500)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_CO5),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_AO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.I5(CLBLM_R_X7Y149_SLICE_X8Y149_CO6),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303003301010011)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd4dc777fd7df575f)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h080000ccf000f000)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3322110033321110)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_DO6),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_AO5),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_BO6),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_BO5),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_BO5),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_AO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfff4fffcffe4ffe)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbf4f8f3fff0fcf)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_DO6),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7757ff33775733ff)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_BLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.I1(CLBLM_R_X7Y150_SLICE_X9Y150_BO6),
.I2(CLBLM_L_X16Y142_SLICE_X22Y142_AO5),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccfffccccffff)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_CO6),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_BO6),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I5(CLBLM_R_X7Y150_SLICE_X8Y150_CO6),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_AO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3323333333013331)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffcaff8f)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_CLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888800005555)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f0eefffeff)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_CO6),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8844fffff0f0ffff)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_CO5),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_BO6),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000022aa000033f3)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500af0005050505)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h222e222e222e000c)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_DO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I3(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_CO6),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcacdcfcdc)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_CO5),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.I4(CLBLM_R_X7Y151_SLICE_X8Y151_BO5),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y130_SLICE_X14Y130_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X11Y130_SLICE_X14Y130_D_CY, CLBLM_R_X11Y130_SLICE_X14Y130_C_CY, CLBLM_R_X11Y130_SLICE_X14Y130_B_CY, CLBLM_R_X11Y130_SLICE_X14Y130_A_CY}),
.CYINIT(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.DI({1'b0, 1'b0, 1'b0, CLBLM_R_X11Y130_SLICE_X14Y130_AO5}),
.O({CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR, CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR, CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR, CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR}),
.S({CLBLM_R_X11Y130_SLICE_X14Y130_DO6, CLBLM_R_X11Y130_SLICE_X14Y130_CO6, CLBLM_R_X11Y130_SLICE_X14Y130_BO6, CLBLM_R_X11Y130_SLICE_X14Y130_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y130_SLICE_X15Y130_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X11Y130_SLICE_X15Y130_D_CY, CLBLM_R_X11Y130_SLICE_X15Y130_C_CY, CLBLM_R_X11Y130_SLICE_X15Y130_B_CY, CLBLM_R_X11Y130_SLICE_X15Y130_A_CY}),
.CYINIT(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.DI({1'b0, 1'b0, 1'b0, CLBLM_R_X11Y130_SLICE_X15Y130_AO5}),
.O({CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR, CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR, CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR, CLBLM_R_X11Y130_SLICE_X15Y130_A_XOR}),
.S({CLBLM_R_X11Y130_SLICE_X15Y130_DO6, CLBLM_R_X11Y130_SLICE_X15Y130_CO6, CLBLM_R_X11Y130_SLICE_X15Y130_BO6, CLBLM_R_X11Y130_SLICE_X15Y130_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_BQ),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CARRY4 (
.CI(CLBLM_R_X11Y130_SLICE_X14Y130_COUT),
.CO({CLBLM_R_X11Y131_SLICE_X14Y131_D_CY, CLBLM_R_X11Y131_SLICE_X14Y131_C_CY, CLBLM_R_X11Y131_SLICE_X14Y131_B_CY, CLBLM_R_X11Y131_SLICE_X14Y131_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR, CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR, CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR, CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR}),
.S({CLBLM_R_X11Y131_SLICE_X14Y131_DO6, CLBLM_R_X11Y131_SLICE_X14Y131_CO6, CLBLM_R_X11Y131_SLICE_X14Y131_BO6, CLBLM_R_X11Y131_SLICE_X14Y131_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CARRY4 (
.CI(CLBLM_R_X11Y130_SLICE_X15Y130_COUT),
.CO({CLBLM_R_X11Y131_SLICE_X15Y131_D_CY, CLBLM_R_X11Y131_SLICE_X15Y131_C_CY, CLBLM_R_X11Y131_SLICE_X15Y131_B_CY, CLBLM_R_X11Y131_SLICE_X15Y131_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR, CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR, CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR, CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR}),
.S({CLBLM_R_X11Y131_SLICE_X15Y131_DO6, CLBLM_R_X11Y131_SLICE_X15Y131_CO6, CLBLM_R_X11Y131_SLICE_X15Y131_BO6, CLBLM_R_X11Y131_SLICE_X15Y131_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_A5Q),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y132_SLICE_X14Y132_AO5),
.Q(CLBLM_R_X11Y132_SLICE_X14Y132_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y132_SLICE_X14Y132_CARRY4 (
.CI(CLBLM_R_X11Y131_SLICE_X14Y131_COUT),
.CO({CLBLM_R_X11Y132_SLICE_X14Y132_D_CY, CLBLM_R_X11Y132_SLICE_X14Y132_C_CY, CLBLM_R_X11Y132_SLICE_X14Y132_B_CY, CLBLM_R_X11Y132_SLICE_X14Y132_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR, CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR, CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR, CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR}),
.S({CLBLM_R_X11Y132_SLICE_X14Y132_DO6, CLBLM_R_X11Y132_SLICE_X14Y132_CO6, CLBLM_R_X11Y132_SLICE_X14Y132_BO6, CLBLM_R_X11Y132_SLICE_X14Y132_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_A5Q),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_A5Q),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y132_SLICE_X15Y132_CARRY4 (
.CI(CLBLM_R_X11Y131_SLICE_X15Y131_COUT),
.CO({CLBLM_R_X11Y132_SLICE_X15Y132_D_CY, CLBLM_R_X11Y132_SLICE_X15Y132_C_CY, CLBLM_R_X11Y132_SLICE_X15Y132_B_CY, CLBLM_R_X11Y132_SLICE_X15Y132_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR, CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR, CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR, CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR}),
.S({CLBLM_R_X11Y132_SLICE_X15Y132_DO6, CLBLM_R_X11Y132_SLICE_X15Y132_CO6, CLBLM_R_X11Y132_SLICE_X15Y132_BO6, CLBLM_R_X11Y132_SLICE_X15Y132_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_A5Q),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_B5Q),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y131_SLICE_X17Y131_A5Q),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y133_SLICE_X14Y133_CARRY4 (
.CI(CLBLM_R_X11Y132_SLICE_X14Y132_COUT),
.CO({CLBLM_R_X11Y133_SLICE_X14Y133_D_CY, CLBLM_R_X11Y133_SLICE_X14Y133_C_CY, CLBLM_R_X11Y133_SLICE_X14Y133_B_CY, CLBLM_R_X11Y133_SLICE_X14Y133_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y133_SLICE_X14Y133_D_XOR, CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR, CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR, CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR}),
.S({CLBLM_R_X11Y133_SLICE_X14Y133_DO6, CLBLM_R_X11Y133_SLICE_X14Y133_CO6, CLBLM_R_X11Y133_SLICE_X14Y133_BO6, CLBLM_R_X11Y133_SLICE_X14Y133_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y131_SLICE_X16Y131_A5Q),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_B5Q),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y132_SLICE_X17Y132_BQ),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y133_SLICE_X15Y133_CARRY4 (
.CI(CLBLM_R_X11Y132_SLICE_X15Y132_COUT),
.CO({CLBLM_R_X11Y133_SLICE_X15Y133_D_CY, CLBLM_R_X11Y133_SLICE_X15Y133_C_CY, CLBLM_R_X11Y133_SLICE_X15Y133_B_CY, CLBLM_R_X11Y133_SLICE_X15Y133_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y133_SLICE_X15Y133_D_XOR, CLBLM_R_X11Y133_SLICE_X15Y133_C_XOR, CLBLM_R_X11Y133_SLICE_X15Y133_B_XOR, CLBLM_R_X11Y133_SLICE_X15Y133_A_XOR}),
.S({CLBLM_R_X11Y133_SLICE_X15Y133_DO6, CLBLM_R_X11Y133_SLICE_X15Y133_CO6, CLBLM_R_X11Y133_SLICE_X15Y133_BO6, CLBLM_R_X11Y133_SLICE_X15Y133_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0035f0350f35ff35)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_DLUT (
.I0(CLBLL_L_X26Y133_SLICE_X38Y133_CO5),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h353500f035350fff)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_CLUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I5(CLBLL_L_X26Y133_SLICE_X38Y133_CO6),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e2e2f0f0f0aa)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_BLUT (
.I0(CLBLL_L_X26Y133_SLICE_X38Y133_BO5),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I2(CLBLL_L_X26Y133_SLICE_X38Y133_BO6),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff02fd00ff07f800)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I3(CLBLL_L_X26Y133_SLICE_X38Y133_CO6),
.I4(CLBLL_L_X26Y133_SLICE_X38Y133_CO5),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.Q(CLBLM_R_X11Y134_SLICE_X15Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333f0aaf000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_DLUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_AQ),
.I1(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_CO6),
.I4(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccaa00f0ccaaff)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_CLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_AO6),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_BO6),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_DO6),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0b8f0f0e2aa)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_BLUT (
.I0(CLBLL_L_X26Y133_SLICE_X38Y133_DO5),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I2(CLBLL_L_X26Y133_SLICE_X38Y133_DO6),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000fffffb8b8b8b8)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_ALUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_DO6),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_CO6),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I3(CLBLM_R_X11Y135_SLICE_X15Y135_CQ),
.I4(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y135_SLICE_X14Y135_AO6),
.Q(CLBLM_R_X11Y135_SLICE_X14Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccf0f05555)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_DLUT (
.I0(CLBLM_R_X11Y135_SLICE_X15Y135_CQ),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_CO6),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_AO5),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_DO6),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefab6723cd894501)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_BO6),
.I4(CLBLM_R_X7Y135_SLICE_X8Y135_BO6),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_BO6),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c11dd3f3f11dd)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_BLUT (
.I0(CLBLL_L_X26Y133_SLICE_X38Y133_AO5),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I5(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf030f0b8f0fcf0b8)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_AO6),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y135_SLICE_X15Y135_BO6),
.Q(CLBLM_R_X11Y135_SLICE_X15Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y135_SLICE_X15Y135_CO6),
.Q(CLBLM_R_X11Y135_SLICE_X15Y135_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0aaccaacc)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_DLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I2(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I4(CLBLM_R_X11Y135_SLICE_X15Y135_CQ),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0acc0fccfaccffcc)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X11Y135_SLICE_X15Y135_CQ),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_DO6),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_CO6),
.I5(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ee44cccc)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_BLUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I1(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_DO6),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c3f0c3faaaaeeee)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_ALUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_A5Q),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.Q(CLBLM_R_X11Y136_SLICE_X14Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y136_SLICE_X14Y136_BO6),
.Q(CLBLM_R_X11Y136_SLICE_X14Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f3fffff7733ffff)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f1e0f0f0fd20)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_CLUT (
.I0(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I2(CLBLL_L_X26Y133_SLICE_X38Y133_AO6),
.I3(CLBLL_L_X26Y133_SLICE_X38Y133_AO5),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddd8d8d8d8)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.I1(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.I2(CLBLM_R_X11Y136_SLICE_X15Y136_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y135_SLICE_X8Y135_CO6),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8bbb8bbb888b888)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_ALUT (
.I0(CLBLM_L_X12Y146_SLICE_X17Y146_CO6),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.I2(CLBLM_R_X13Y136_SLICE_X18Y136_DO6),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AO5),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y136_SLICE_X15Y136_AO6),
.Q(CLBLM_R_X11Y136_SLICE_X15Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y136_SLICE_X15Y136_BO6),
.Q(CLBLM_R_X11Y136_SLICE_X15Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb000000000000000)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002070f0f02070)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_CLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_DO6),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_DO6),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I5(CLBLM_R_X13Y135_SLICE_X18Y135_DO6),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8cdcdcdc8cdc8c8c)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_BLUT (
.I0(CLBLM_L_X12Y137_SLICE_X16Y137_CO6),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I3(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h77f0f0f044f0f0f0)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_ALUT (
.I0(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.I2(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_BO6),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffac0facf0ac00ac)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_DO6),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_CO6),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I4(CLBLM_L_X10Y137_SLICE_X12Y137_DO6),
.I5(CLBLM_R_X7Y137_SLICE_X9Y137_BO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcffa0ac0c0fa0a)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_CLUT (
.I0(CLBLM_R_X11Y137_SLICE_X15Y137_BO6),
.I1(CLBLM_L_X16Y137_SLICE_X22Y137_CO6),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I3(CLBLM_R_X13Y137_SLICE_X18Y137_AO6),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I5(CLBLM_L_X16Y137_SLICE_X22Y137_DO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h048c26ae159d37bf)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_BLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.I2(CLBLM_R_X15Y137_SLICE_X21Y137_CO6),
.I3(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I4(CLBLM_R_X13Y137_SLICE_X18Y137_BO6),
.I5(CLBLM_L_X16Y134_SLICE_X22Y134_CO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a01111bbbb)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_BO6),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X11Y137_SLICE_X14Y137_MUXF7A (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_BO6),
.I1(CLBLM_R_X11Y137_SLICE_X14Y137_AO6),
.O(CLBLM_R_X11Y137_SLICE_X14Y137_F7AMUX_O),
.S(CLBLM_R_X11Y143_SLICE_X14Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_R_X11Y137_SLICE_X14Y137_MUXF7B (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_DO6),
.I1(CLBLM_R_X11Y137_SLICE_X14Y137_CO6),
.O(CLBLM_R_X11Y137_SLICE_X14Y137_F7BMUX_O),
.S(CLBLM_R_X11Y143_SLICE_X14Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_R_X11Y137_SLICE_X14Y137_MUXF8 (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_F7BMUX_O),
.I1(CLBLM_R_X11Y137_SLICE_X14Y137_F7AMUX_O),
.O(CLBLM_R_X11Y137_SLICE_X14Y137_F8MUX_O),
.S(CLBLM_R_X7Y141_SLICE_X8Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff05fa00ff03fc00)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I1(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_AO6),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd080df8f00000f0f)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I1(CLBLM_R_X11Y135_SLICE_X15Y135_DO6),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.DIB(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.DIC(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.DID(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.DOA(CLBLM_R_X11Y138_SLICE_X14Y138_AO6),
.DOB(CLBLM_R_X11Y138_SLICE_X14Y138_BO6),
.DOC(CLBLM_R_X11Y138_SLICE_X14Y138_CO6),
.DOD(CLBLM_R_X11Y138_SLICE_X14Y138_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_L_X12Y140_SLICE_X17Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y138_SLICE_X15Y138_AO6),
.Q(CLBLM_R_X11Y138_SLICE_X15Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555d1d1d1d1)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_DO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff270027ff270027)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_CLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I2(CLBLM_R_X13Y138_SLICE_X18Y138_DO6),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_CO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff3fff00ff0f)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y138_SLICE_X17Y138_AO6),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_BO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fa50fa50fa50)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_ALUT (
.I0(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.I3(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_DO6),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_AO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.DIB(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.DIC(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.DID(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.DOA(CLBLM_R_X11Y139_SLICE_X14Y139_AO6),
.DOB(CLBLM_R_X11Y139_SLICE_X14Y139_BO6),
.DOC(CLBLM_R_X11Y139_SLICE_X14Y139_CO6),
.DOD(CLBLM_R_X11Y139_SLICE_X14Y139_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_L_X12Y139_SLICE_X17Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y139_SLICE_X15Y139_AO6),
.Q(CLBLM_R_X11Y139_SLICE_X15Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y139_SLICE_X15Y139_BO6),
.Q(CLBLM_R_X11Y139_SLICE_X15Y139_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f5555000f5555)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_DO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_AO6),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_CO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030bb88bb88)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_BLUT (
.I0(CLBLM_L_X12Y138_SLICE_X16Y138_AO6),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_AO6),
.I3(CLBLM_R_X13Y139_SLICE_X18Y139_AO6),
.I4(CLBLM_R_X11Y138_SLICE_X14Y138_AO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_BO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ccaaccaa)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_ALUT (
.I0(CLBLM_R_X13Y139_SLICE_X18Y139_CO6),
.I1(CLBLM_L_X12Y138_SLICE_X16Y138_CO6),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_CO6),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.I4(CLBLM_R_X11Y138_SLICE_X14Y138_CO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_AO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X12Y140_SLICE_X17Y140_CO6),
.DIB(CLBLM_L_X12Y142_SLICE_X17Y142_DO6),
.DIC(CLBLM_R_X13Y141_SLICE_X18Y141_BO6),
.DID(1'b0),
.DOA(CLBLM_R_X11Y140_SLICE_X14Y140_AO6),
.DOB(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.DOC(CLBLM_R_X11Y140_SLICE_X14Y140_CO6),
.DOD(CLBLM_R_X11Y140_SLICE_X14Y140_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_R_X11Y139_SLICE_X15Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_AO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_BO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_CO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_DO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0fff000)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_DLUT (
.I0(CLBLM_L_X12Y140_SLICE_X16Y140_CO6),
.I1(CLBLM_L_X12Y139_SLICE_X16Y139_CO6),
.I2(CLBLM_L_X12Y141_SLICE_X16Y141_CO6),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_CO6),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_DO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33b8b8cc00b8b8)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_CLUT (
.I0(CLBLM_L_X12Y139_SLICE_X16Y139_BO6),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.I2(CLBLM_R_X13Y140_SLICE_X18Y140_BO6),
.I3(CLBLM_L_X12Y140_SLICE_X16Y140_BO6),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I5(CLBLM_L_X12Y141_SLICE_X16Y141_BO6),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_CO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888f3c0f3c0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_BLUT (
.I0(CLBLM_L_X12Y140_SLICE_X16Y140_AO6),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.I2(CLBLM_L_X12Y139_SLICE_X16Y139_AO6),
.I3(CLBLM_R_X13Y140_SLICE_X18Y140_AO6),
.I4(CLBLM_L_X12Y141_SLICE_X16Y141_AO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_BO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88f3f3bb88c0c0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_ALUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_CO6),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_CO6),
.I3(CLBLM_R_X11Y141_SLICE_X14Y141_CO6),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I5(CLBLM_L_X12Y142_SLICE_X16Y142_CO6),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_AO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X12Y140_SLICE_X17Y140_CO6),
.DIB(CLBLM_L_X12Y142_SLICE_X17Y142_DO6),
.DIC(CLBLM_R_X13Y141_SLICE_X18Y141_BO6),
.DID(CLBLM_R_X11Y143_SLICE_X15Y143_DO6),
.DOA(CLBLM_R_X11Y141_SLICE_X14Y141_AO6),
.DOB(CLBLM_R_X11Y141_SLICE_X14Y141_BO6),
.DOC(CLBLM_R_X11Y141_SLICE_X14Y141_CO6),
.DOD(CLBLM_R_X11Y141_SLICE_X14Y141_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_L_X12Y139_SLICE_X17Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y142_SLICE_X18Y142_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0faa0f550f000f)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_DLUT (
.I0(CLBLM_L_X12Y141_SLICE_X17Y141_AO6),
.I1(1'b1),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_BO5),
.I5(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_DO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccf0f0aaaa)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_CLUT (
.I0(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I1(CLBLM_R_X11Y140_SLICE_X15Y140_DQ),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_DQ),
.I3(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_CO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_BLUT (
.I0(CLBLM_R_X11Y143_SLICE_X15Y143_A5Q),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_CQ),
.I4(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_BO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfc0cfc0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_ALUT (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_CQ),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_AO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X12Y140_SLICE_X17Y140_CO6),
.DIB(CLBLM_L_X12Y142_SLICE_X17Y142_DO6),
.DIC(CLBLM_R_X13Y141_SLICE_X18Y141_BO6),
.DID(1'b0),
.DOA(CLBLM_R_X11Y142_SLICE_X14Y142_AO6),
.DOB(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.DOC(CLBLM_R_X11Y142_SLICE_X14Y142_CO6),
.DOD(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_L_X12Y140_SLICE_X17Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y140_SLICE_X17Y140_CO6),
.Q(CLBLM_R_X11Y142_SLICE_X15Y142_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00f0f0aaaa)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I2(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_DO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaccccf0f0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_CLUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_A5Q),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_CO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0bbbbf3c08888)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_BLUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_DQ),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I2(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(CLBLM_R_X11Y140_SLICE_X15Y140_CQ),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_BO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888f3c0f3c0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_ALUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_DQ),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_CQ),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_AO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X11Y142_SLICE_X15Y142_MUXF7A (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_BO6),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_AO6),
.O(CLBLM_R_X11Y142_SLICE_X15Y142_F7AMUX_O),
.S(CLBLM_L_X10Y139_SLICE_X12Y139_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_R_X11Y142_SLICE_X15Y142_MUXF7B (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_DO6),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_CO6),
.O(CLBLM_R_X11Y142_SLICE_X15Y142_F7BMUX_O),
.S(CLBLM_L_X10Y139_SLICE_X12Y139_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_R_X11Y142_SLICE_X15Y142_MUXF8 (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_F7BMUX_O),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_F7AMUX_O),
.O(CLBLM_R_X11Y142_SLICE_X15Y142_F8MUX_O),
.S(CLBLM_R_X11Y141_SLICE_X15Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfccafaac0cca0aa)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_DLUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_A5Q),
.I2(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I3(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(CLBLM_L_X10Y137_SLICE_X13Y137_BQ),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeff4400e4f0e4f0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_CLUT (
.I0(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I1(CLBLM_L_X10Y137_SLICE_X13Y137_CQ),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_DQ),
.I3(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I4(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcb87430ffaa5500)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_BLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_CQ),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I5(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0704f7f4)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_ALUT (
.I0(CLBLM_R_X15Y141_SLICE_X20Y141_DO6),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_AO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y141_SLICE_X18Y141_BO6),
.Q(CLBLM_R_X11Y143_SLICE_X15Y143_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y143_SLICE_X15Y143_AO6),
.Q(CLBLM_R_X11Y143_SLICE_X15Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aafceef0aa3022)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_CLUT (
.I0(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_DQ),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I4(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I5(CLBLM_R_X11Y136_SLICE_X14Y136_BQ),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfd0808fd08fd08)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_BLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.I2(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I3(CLBLM_R_X11Y142_SLICE_X15Y142_F7BMUX_O),
.I4(CLBLM_R_X11Y142_SLICE_X15Y142_F7AMUX_O),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff88000f00)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_CLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I1(CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_AO6),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_BO6),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff2fff2fff20f02)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_BLUT (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_BO6),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AO6),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_BO6),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80808080ffff55ff)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfff2fffffffffff)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_AO6),
.I3(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_BO6),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c000c0044000000)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_CLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f66ffff0f66ff00)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_BLUT (
.I0(CLBLM_R_X11Y145_SLICE_X14Y145_DO6),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_AO6),
.I2(CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccfeeef00032223)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_ALUT (
.I0(CLBLM_L_X12Y147_SLICE_X16Y147_BQ),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_BO6),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_BO5),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_CO6),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecccefccdcccdfcc)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_BLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_CO6),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_CO6),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I3(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I5(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf773000031100000)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_AO6),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c555caaacfff)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR),
.I5(CLBLM_R_X13Y146_SLICE_X18Y146_C_XOR),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ccc0c440c880c00)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I4(CLBLM_R_X13Y146_SLICE_X18Y146_B_XOR),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fcf0fc000c505c)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_BLUT (
.I0(CLBLM_R_X15Y149_SLICE_X20Y149_AO5),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_BO5),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_CO6),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8083b0b300000000)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_ALUT (
.I0(CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_AO6),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdef05af012305af)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR),
.I3(CLBLM_R_X13Y146_SLICE_X18Y146_A_XOR),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a022772277)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_R_X13Y146_SLICE_X18Y146_D_XOR),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeeef0f0fff0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_BLUT (
.I0(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_AO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00110001)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_ALUT (
.I0(CLBLM_R_X13Y147_SLICE_X19Y147_CO6),
.I1(CLBLM_R_X13Y148_SLICE_X18Y148_BO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I4(CLBLM_R_X13Y146_SLICE_X19Y146_BO6),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h555555550f0f0f0f)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfff0aacc00f0aa)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I2(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacac00f0acac0fff)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I3(CLBLM_R_X13Y147_SLICE_X18Y147_A_XOR),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800f7ff8c0073ff)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_ALUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I1(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_BO6),
.I4(CLBLM_R_X7Y145_SLICE_X9Y145_AO6),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_DQ),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80007f004000bf00)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_DLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I5(CLBLM_R_X11Y150_SLICE_X14Y150_AO5),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff888888fff8f8f8)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_CLUT (
.I0(CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I3(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I4(CLBLM_R_X13Y146_SLICE_X19Y146_AO5),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_BO6),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdf0fdfffffffff)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_CO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa0eca0eca0ec)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_ALUT (
.I0(CLBLM_L_X12Y147_SLICE_X16Y147_CQ),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I2(CLBLM_R_X13Y146_SLICE_X19Y146_AO5),
.I3(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.I4(CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000c400000080)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_DLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_BO6),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fff3ffbbffffff)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb24d4db24dff004d)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_BLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c080808080)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_CQ),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0000020200000)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_DLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_DO6),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeac0ffffc0c0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_CLUT (
.I0(CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR),
.I1(CLBLM_R_X13Y146_SLICE_X19Y146_AO5),
.I2(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.I4(CLBLM_R_X11Y148_SLICE_X15Y148_DO6),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_AO5),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeac0c0ffeaffc0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_BLUT (
.I0(CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR),
.I1(CLBLM_R_X13Y146_SLICE_X19Y146_AO5),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_BO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeeafaacfcc0f00)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_ALUT (
.I0(CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR),
.I1(CLBLM_R_X13Y146_SLICE_X19Y146_AO5),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_CO6),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_DQ),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_CO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_DO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b4f0f0f0f0f0f0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_DLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc9ccccccccccccc)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c33c698e0ccf8e)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_BLUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc006c9336c9)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0afa0ff00ff00)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_DLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_BO6),
.I1(CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_DO6),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaacd5522aa0155)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h300a3f0a30fa3ffa)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(CLBLM_L_X12Y144_SLICE_X17Y144_DO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_BO6),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_CO6),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800240000000800)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdfdf8080dfdfdf)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_DO6),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_AO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fe070effff0f0f)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_CLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I4(CLBLM_R_X11Y150_SLICE_X14Y150_DO6),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0517175f71f55071)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h872d0f0f3f033f03)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c3693c933333333)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_DLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9555a9999995aaa9)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_CLUT (
.I0(CLBLM_R_X11Y150_SLICE_X15Y150_AO6),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5f54050fdff5455)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I1(CLBLM_R_X11Y145_SLICE_X15Y145_AO6),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I3(CLBLM_R_X15Y151_SLICE_X20Y151_AO6),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff00054d4d5f)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_AO5),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_BO5),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_AO6),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y128_SLICE_X18Y128_BO6),
.Q(CLBLM_R_X13Y128_SLICE_X18Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000002)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_CLUT (
.I0(CLBLM_L_X12Y129_SLICE_X17Y129_AO6),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I3(CLBLM_R_X13Y128_SLICE_X18Y128_A5Q),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h003c00cc006a00aa)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_BLUT (
.I0(CLBLM_R_X13Y128_SLICE_X18Y128_B5Q),
.I1(CLBLM_R_X13Y128_SLICE_X18Y128_BQ),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050505055050)
  ) CLBLM_R_X13Y128_SLICE_X18Y128_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I1(1'b1),
.I2(CLBLM_R_X13Y128_SLICE_X18Y128_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y128_SLICE_X18Y128_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X18Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X18Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_DO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_CO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_BO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y128_SLICE_X19Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y128_SLICE_X19Y128_AO5),
.O6(CLBLM_R_X13Y128_SLICE_X19Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y129_SLICE_X18Y129_BO5),
.Q(CLBLM_R_X13Y129_SLICE_X18Y129_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y129_SLICE_X18Y129_AO6),
.Q(CLBLM_R_X13Y129_SLICE_X18Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y129_SLICE_X18Y129_BO6),
.Q(CLBLM_R_X13Y129_SLICE_X18Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y129_SLICE_X18Y129_CO6),
.Q(CLBLM_R_X13Y129_SLICE_X18Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000000080000)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I3(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6060c0c0c0c0c0c0)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_CLUT (
.I0(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_CQ),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I3(1'b1),
.I4(CLBLM_R_X13Y129_SLICE_X18Y129_B5Q),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3330000066600000)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_BLUT (
.I0(CLBLM_R_X13Y129_SLICE_X18Y129_B5Q),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0078000000780000)
  ) CLBLM_R_X13Y129_SLICE_X18Y129_ALUT (
.I0(CLBLM_R_X13Y129_SLICE_X18Y129_B5Q),
.I1(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I2(CLBLM_R_X13Y129_SLICE_X18Y129_AQ),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_BO6),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X18Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X18Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y129_SLICE_X19Y129_AO6),
.Q(CLBLM_R_X13Y129_SLICE_X19Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a08080a0a08080)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_DLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_DO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fca80000)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_CLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I3(CLBLM_R_X13Y136_SLICE_X19Y136_BQ),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I5(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_CO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f4f5f7f00300000)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_BLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_BO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000c0000000c)
  ) CLBLM_R_X13Y129_SLICE_X19Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y130_SLICE_X18Y130_BO6),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I3(CLBLM_R_X13Y129_SLICE_X19Y129_BO6),
.I4(CLBLM_R_X15Y129_SLICE_X20Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y129_SLICE_X19Y129_AO5),
.O6(CLBLM_R_X13Y129_SLICE_X19Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y130_SLICE_X18Y130_AO6),
.Q(CLBLM_R_X13Y130_SLICE_X18Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5554545454545454)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_DLUT (
.I0(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I1(CLBLM_R_X13Y130_SLICE_X19Y130_CO6),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_BO5),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_CQ),
.I4(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I5(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050000000400000)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_CLUT (
.I0(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_CQ),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef4fcfcf4f4fcfc)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_BLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I1(CLBLM_R_X13Y136_SLICE_X19Y136_BQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_BO6),
.I3(CLBLM_R_X13Y129_SLICE_X18Y129_BQ),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I5(CLBLM_R_X13Y129_SLICE_X18Y129_CQ),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaf000faaa0000)
  ) CLBLM_R_X13Y130_SLICE_X18Y130_ALUT (
.I0(CLBLM_R_X13Y129_SLICE_X19Y129_BO5),
.I1(1'b1),
.I2(CLBLM_L_X12Y129_SLICE_X17Y129_AQ),
.I3(CLBLM_R_X13Y129_SLICE_X19Y129_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_L_X12Y130_SLICE_X17Y130_AQ),
.O5(CLBLM_R_X13Y130_SLICE_X18Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X18Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y130_SLICE_X19Y130_AO6),
.Q(CLBLM_R_X13Y130_SLICE_X19Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_DO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0d100000000)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_CLUT (
.I0(CLBLM_L_X16Y136_SLICE_X22Y136_BQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I5(CLBLM_R_X13Y136_SLICE_X19Y136_BQ),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_CO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfffdffa8aafdff)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_BLUT (
.I0(CLBLM_R_X15Y131_SLICE_X21Y131_BO6),
.I1(CLBLM_L_X16Y136_SLICE_X22Y136_BQ),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I3(CLBLM_R_X13Y136_SLICE_X19Y136_BQ),
.I4(CLBLM_R_X15Y130_SLICE_X20Y130_AQ),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_BO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ff0000f0f0)
  ) CLBLM_R_X13Y130_SLICE_X19Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I3(CLBLM_R_X13Y130_SLICE_X19Y130_BO6),
.I4(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_CO6),
.O5(CLBLM_R_X13Y130_SLICE_X19Y130_AO5),
.O6(CLBLM_R_X13Y130_SLICE_X19Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y131_SLICE_X20Y131_AQ),
.Q(CLBLM_R_X13Y131_SLICE_X18Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y131_SLICE_X19Y131_BQ),
.Q(CLBLM_R_X13Y131_SLICE_X18Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y131_SLICE_X19Y131_DQ),
.Q(CLBLM_R_X13Y131_SLICE_X18Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.Q(CLBLM_R_X13Y131_SLICE_X18Y131_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_DO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800000000000)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_CO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffbfffffffffff)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_BLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_A5Q),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y130_SLICE_X16Y130_CQ),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_BO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11cc44f0f0f0f0)
  ) CLBLM_R_X13Y131_SLICE_X18Y131_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X17Y131_DO6),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR),
.I3(CLBLM_R_X13Y131_SLICE_X18Y131_BO6),
.I4(CLBLM_R_X13Y131_SLICE_X18Y131_CO6),
.I5(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.O5(CLBLM_R_X13Y131_SLICE_X18Y131_AO5),
.O6(CLBLM_R_X13Y131_SLICE_X18Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y131_SLICE_X19Y131_AO6),
.Q(CLBLM_R_X13Y131_SLICE_X19Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y131_SLICE_X19Y131_BO6),
.Q(CLBLM_R_X13Y131_SLICE_X19Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y131_SLICE_X19Y131_CO6),
.Q(CLBLM_R_X13Y131_SLICE_X19Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y131_SLICE_X19Y131_DO6),
.Q(CLBLM_R_X13Y131_SLICE_X19Y131_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc000400c8000000)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_DLUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I1(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_AQ),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I5(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_DO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32fefafa32fafa)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_CLUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I1(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I3(CLBLM_R_X13Y131_SLICE_X19Y131_DQ),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I5(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_CO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f3ffffffff)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_BLUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I2(CLBLM_R_X13Y131_SLICE_X19Y131_CQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I5(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_BO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888c000088800000)
  ) CLBLM_R_X13Y131_SLICE_X19Y131_ALUT (
.I0(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I1(CLBLM_R_X13Y130_SLICE_X18Y130_AQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I5(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.O5(CLBLM_R_X13Y131_SLICE_X19Y131_AO5),
.O6(CLBLM_R_X13Y131_SLICE_X19Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y132_SLICE_X18Y132_DO5),
.Q(CLBLM_R_X13Y132_SLICE_X18Y132_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y132_SLICE_X18Y132_DO6),
.Q(CLBLM_R_X13Y132_SLICE_X18Y132_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333030fcfc0303)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y133_SLICE_X17Y133_CO6),
.I2(CLBLM_R_X13Y135_SLICE_X19Y135_DQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfc0cfc0)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_CLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_L_X12Y131_SLICE_X17Y131_A5Q),
.I4(CLBLM_L_X12Y132_SLICE_X17Y132_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h330033ffaaf0aaf0)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I1(CLBLM_R_X13Y138_SLICE_X18Y138_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X17Y131_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I4(CLBLM_R_X13Y134_SLICE_X19Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0cc00cc00)
  ) CLBLM_R_X13Y132_SLICE_X18Y132_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I3(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X18Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X18Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_DO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_CO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_BO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y132_SLICE_X19Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y132_SLICE_X19Y132_AO5),
.O6(CLBLM_R_X13Y132_SLICE_X19Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_DO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22f3f3ee22c0c0)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_CLUT (
.I0(CLBLM_R_X15Y134_SLICE_X21Y134_BQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_CO6),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.I5(CLBLM_R_X15Y136_SLICE_X21Y136_CQ),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_CO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h53535353000ff0ff)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_BLUT (
.I0(CLBLM_R_X13Y136_SLICE_X18Y136_B5Q),
.I1(CLBLM_R_X13Y133_SLICE_X19Y133_B5Q),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X13Y134_SLICE_X19Y134_BQ),
.I4(CLBLM_L_X12Y138_SLICE_X17Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_BO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc33ffe2e2e2e2)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_ALUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_AQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I3(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.I4(CLBLM_R_X13Y133_SLICE_X19Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_AO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y133_SLICE_X19Y133_AO5),
.Q(CLBLM_R_X13Y133_SLICE_X19Y133_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y133_SLICE_X19Y133_BO5),
.Q(CLBLM_R_X13Y133_SLICE_X19Y133_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y133_SLICE_X19Y133_AO6),
.Q(CLBLM_R_X13Y133_SLICE_X19Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y133_SLICE_X19Y133_BO6),
.Q(CLBLM_R_X13Y133_SLICE_X19Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00110005eefffaff)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_DLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I2(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I3(CLBLM_R_X13Y136_SLICE_X19Y136_AQ),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I5(CLBLM_L_X16Y136_SLICE_X23Y136_AQ),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_DO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f0f0f0000)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.I3(1'b1),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4e4e4e4e55ff00aa)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.I1(CLBLM_R_X15Y133_SLICE_X21Y133_BQ),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I4(CLBLM_R_X15Y133_SLICE_X21Y133_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_BO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dd88dd88)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.I1(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I3(CLBLM_R_X15Y134_SLICE_X21Y134_BQ),
.I4(CLBLM_R_X15Y133_SLICE_X21Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_AO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333001033330000)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_DLUT (
.I0(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_DO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccdccccccccc)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_CO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333ccceccce)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_BLUT (
.I0(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I1(CLBLM_R_X13Y134_SLICE_X19Y134_DO6),
.I2(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I4(CLBLM_R_X15Y137_SLICE_X20Y137_D_CY),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f00fff35353535)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_ALUT (
.I0(CLBLM_R_X13Y133_SLICE_X19Y133_A5Q),
.I1(CLBLM_R_X13Y136_SLICE_X18Y136_A5Q),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_R_X13Y136_SLICE_X18Y136_BQ),
.I4(CLBLM_R_X13Y133_SLICE_X19Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_AO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y134_SLICE_X19Y134_AO5),
.Q(CLBLM_R_X13Y134_SLICE_X19Y134_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y134_SLICE_X19Y134_BO5),
.Q(CLBLM_R_X13Y134_SLICE_X19Y134_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y134_SLICE_X19Y134_AO6),
.Q(CLBLM_R_X13Y134_SLICE_X19Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y134_SLICE_X19Y134_BO6),
.Q(CLBLM_R_X13Y134_SLICE_X19Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7ffffffffff)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_DLUT (
.I0(CLBLM_R_X15Y133_SLICE_X21Y133_BQ),
.I1(CLBLM_R_X15Y136_SLICE_X21Y136_BQ),
.I2(CLBLM_R_X15Y135_SLICE_X21Y135_CO6),
.I3(CLBLM_R_X15Y135_SLICE_X21Y135_BQ),
.I4(CLBLM_R_X13Y135_SLICE_X19Y135_DO6),
.I5(CLBLM_R_X15Y133_SLICE_X21Y133_CQ),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_DO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccaaaaff00)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_CLUT (
.I0(CLBLM_R_X15Y133_SLICE_X21Y133_BQ),
.I1(CLBLM_R_X13Y135_SLICE_X19Y135_CQ),
.I2(CLBLM_R_X13Y132_SLICE_X18Y132_BO5),
.I3(CLBLM_R_X15Y136_SLICE_X21Y136_BQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_CO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222eeee3f0c3f0c)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_BLUT (
.I0(CLBLM_R_X15Y134_SLICE_X21Y134_CQ),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I3(CLBLM_R_X15Y135_SLICE_X21Y135_AQ),
.I4(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_BO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33000faa0faa)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_ALUT (
.I0(CLBLM_R_X15Y135_SLICE_X21Y135_BQ),
.I1(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.I4(CLBLM_R_X15Y134_SLICE_X21Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_AO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.Q(CLBLM_R_X13Y135_SLICE_X18Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_R_X13Y135_SLICE_X18Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80b08cbc83b38fbf)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_DLUT (
.I0(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.I3(CLBLM_R_X15Y135_SLICE_X21Y135_BQ),
.I4(CLBLM_R_X13Y135_SLICE_X19Y135_DQ),
.I5(CLBLM_R_X15Y138_SLICE_X21Y138_BQ),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_DO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222cf03cf03)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_CLUT (
.I0(CLBLM_R_X13Y133_SLICE_X18Y133_AO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_CO6),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_CO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0d1e2e2e2f3)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_BLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I2(CLBLM_R_X13Y135_SLICE_X19Y135_AO6),
.I3(CLBLM_L_X16Y135_SLICE_X22Y135_CO6),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I5(CLBLM_R_X13Y135_SLICE_X18Y135_CO6),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_BO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f00fff53535353)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_ALUT (
.I0(CLBLM_R_X13Y138_SLICE_X18Y138_A5Q),
.I1(CLBLM_R_X13Y134_SLICE_X19Y134_A5Q),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.I3(CLBLM_L_X12Y138_SLICE_X17Y138_BQ),
.I4(CLBLM_R_X13Y134_SLICE_X19Y134_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_AO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.Q(CLBLM_R_X13Y135_SLICE_X19Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.Q(CLBLM_R_X13Y135_SLICE_X19Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_R_X13Y135_SLICE_X19Y135_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_R_X13Y135_SLICE_X19Y135_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffff7f7fffff)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_DLUT (
.I0(CLBLM_R_X15Y133_SLICE_X21Y133_AQ),
.I1(CLBLM_R_X15Y134_SLICE_X21Y134_CQ),
.I2(CLBLM_R_X15Y137_SLICE_X21Y137_AQ),
.I3(1'b1),
.I4(CLBLM_R_X15Y138_SLICE_X21Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_DO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h02075257a2a7f2f7)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.I1(CLBLM_R_X13Y136_SLICE_X19Y136_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.I3(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.I4(CLBLM_R_X15Y134_SLICE_X20Y134_DQ),
.I5(CLBLL_L_X26Y135_SLICE_X38Y135_AO5),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_CO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe5eae04f454a40)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_BLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.I1(CLBLM_R_X13Y135_SLICE_X19Y135_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I3(CLBLM_R_X15Y134_SLICE_X21Y134_AQ),
.I4(CLBLM_R_X15Y137_SLICE_X21Y137_AQ),
.I5(CLBLM_R_X13Y133_SLICE_X18Y133_AO5),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_BO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44ee44)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_ALUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.I1(CLBLM_R_X15Y136_SLICE_X21Y136_AQ),
.I2(CLBLM_R_X13Y135_SLICE_X19Y135_AQ),
.I3(CLBLM_R_X15Y133_SLICE_X21Y133_AQ),
.I4(CLBLM_R_X13Y132_SLICE_X18Y132_AO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_AO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y136_SLICE_X18Y136_AO5),
.Q(CLBLM_R_X13Y136_SLICE_X18Y136_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y136_SLICE_X18Y136_BO5),
.Q(CLBLM_R_X13Y136_SLICE_X18Y136_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y136_SLICE_X18Y136_AO6),
.Q(CLBLM_R_X13Y136_SLICE_X18Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y136_SLICE_X18Y136_BO6),
.Q(CLBLM_R_X13Y136_SLICE_X18Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff001b1b1b1b)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(CLBLM_R_X13Y138_SLICE_X18Y138_CO6),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_BO6),
.I3(CLBLM_R_X13Y136_SLICE_X18Y136_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_DO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef2cec23e320e02)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_CLUT (
.I0(CLBLM_R_X15Y136_SLICE_X21Y136_DQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.I3(CLBLM_R_X15Y133_SLICE_X21Y133_CQ),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_CO5),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_CO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0f0033aa33aa)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_BLUT (
.I0(CLBLM_R_X15Y136_SLICE_X21Y136_DQ),
.I1(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.I4(CLBLM_R_X15Y136_SLICE_X21Y136_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_BO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaa00aa)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_ALUT (
.I0(CLBLM_R_X15Y136_SLICE_X21Y136_CQ),
.I1(CLBLM_R_X15Y136_SLICE_X21Y136_AQ),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_AO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y136_SLICE_X19Y136_AO6),
.Q(CLBLM_R_X13Y136_SLICE_X19Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y136_SLICE_X19Y136_BO6),
.Q(CLBLM_R_X13Y136_SLICE_X19Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaa00aa30)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_BO6),
.I2(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I3(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I4(CLBLM_L_X12Y129_SLICE_X16Y129_BQ),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_DO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fe01ff00ba45ff)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_CLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I2(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I3(CLBLM_R_X13Y136_SLICE_X19Y136_BQ),
.I4(CLBLM_R_X13Y137_SLICE_X19Y137_BQ),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_CO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555fc0c5555cccc)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_BLUT (
.I0(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I1(CLBLM_R_X13Y136_SLICE_X19Y136_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_AO5),
.I3(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I5(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_BO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0aaf0aaf0aa)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_ALUT (
.I0(CLBLM_R_X13Y136_SLICE_X19Y136_AQ),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I4(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.I5(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_AO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y131_SLICE_X19Y131_CQ),
.Q(CLBLM_R_X13Y137_SLICE_X18Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0aff5f000a005f)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y134_SLICE_X17Y134_BO6),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I4(CLBLM_R_X15Y137_SLICE_X21Y137_DO6),
.I5(CLBLM_R_X13Y134_SLICE_X19Y134_CO6),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_DO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500330f55ff330f)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_CLUT (
.I0(CLBLL_L_X26Y136_SLICE_X38Y136_BO5),
.I1(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_BQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.I5(CLBLM_R_X13Y137_SLICE_X19Y137_BQ),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_CO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e2e2f0e2f0e2)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_BLUT (
.I0(CLBLL_L_X26Y136_SLICE_X38Y136_BO5),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLL_L_X26Y136_SLICE_X38Y136_BO6),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_BO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaab8aaaab8b8b8)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_ALUT (
.I0(CLBLL_L_X26Y136_SLICE_X38Y136_AO6),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I2(CLBLM_R_X13Y137_SLICE_X19Y137_AO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_AO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y137_SLICE_X19Y137_BO6),
.Q(CLBLM_R_X13Y137_SLICE_X19Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_DO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_CO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0afa0cfc0cfc0cfc)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_BLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X13Y137_SLICE_X19Y137_BQ),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I3(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.I5(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_BO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505f5f5fe32ce02)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_ALUT (
.I0(CLBLM_R_X13Y138_SLICE_X19Y138_CQ),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_CQ),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_AO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y138_SLICE_X18Y138_AO5),
.Q(CLBLM_R_X13Y138_SLICE_X18Y138_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y138_SLICE_X18Y138_AO6),
.Q(CLBLM_R_X13Y138_SLICE_X18Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0350035ff350f35f)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_DLUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I1(CLBLM_R_X13Y131_SLICE_X18Y131_CQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.I5(CLBLL_L_X26Y138_SLICE_X38Y138_AO6),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_DO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03cf111103cfdddd)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_CLUT (
.I0(CLBLM_L_X12Y137_SLICE_X17Y137_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.I2(CLBLM_R_X13Y136_SLICE_X19Y136_BQ),
.I3(CLBLL_L_X26Y136_SLICE_X38Y136_BO6),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.I5(CLBLM_R_X13Y131_SLICE_X18Y131_BQ),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_CO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e2e2f0f0f0aa)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_BLUT (
.I0(CLBLL_L_X26Y138_SLICE_X38Y138_AO5),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I2(CLBLL_L_X26Y138_SLICE_X38Y138_AO6),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_BO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333f0f05555ff00)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_ALUT (
.I0(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I1(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I2(CLBLM_R_X15Y137_SLICE_X21Y137_AQ),
.I3(CLBLM_R_X15Y138_SLICE_X21Y138_BQ),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_AO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y138_SLICE_X19Y138_AO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X13Y138_SLICE_X19Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_B_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y138_SLICE_X19Y138_BO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X13Y138_SLICE_X19Y138_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_C_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y138_SLICE_X19Y138_CO6),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X13Y138_SLICE_X19Y138_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcfcfcfcfc)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_DO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0cacfcccccccc)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X13Y138_SLICE_X19Y138_CQ),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_DO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_CO6),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_CO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ccd8cc88ccddcc)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.I1(CLBLM_R_X13Y138_SLICE_X19Y138_BQ),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.I4(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_BO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8aaaabb88aaaa)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_ALUT (
.I0(CLBLM_R_X13Y138_SLICE_X19Y138_AQ),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_CO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_AO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.DIB(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.DIC(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.DID(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.DOA(CLBLM_R_X13Y139_SLICE_X18Y139_AO6),
.DOB(CLBLM_R_X13Y139_SLICE_X18Y139_BO6),
.DOC(CLBLM_R_X13Y139_SLICE_X18Y139_CO6),
.DOD(CLBLM_R_X13Y139_SLICE_X18Y139_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_L_X12Y139_SLICE_X17Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e2f0f0f0e2f0)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_DLUT (
.I0(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I1(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I2(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_DO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeedfddeeeedcdd)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_CLUT (
.I0(CLBLM_L_X12Y137_SLICE_X17Y137_AQ),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I5(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_CO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffd)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_BLUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I1(CLBLM_R_X13Y140_SLICE_X19Y140_BO5),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_AO6),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_AO5),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I5(CLBLM_R_X13Y139_SLICE_X19Y139_CO6),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_BO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff1f0e0f0f)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I1(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_AQ),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_AO6)
  );


  (* KEEP, DONT_TOUCH *)
  RAM64M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_RAM64M (
.ADDRA({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRB({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRC({CLBLM_L_X8Y140_SLICE_X10Y140_CO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO6, CLBLM_L_X8Y138_SLICE_X10Y138_DO6, CLBLM_L_X8Y141_SLICE_X11Y141_DO6, CLBLM_L_X10Y141_SLICE_X13Y141_DO6, CLBLM_L_X8Y140_SLICE_X10Y140_DO5}),
.ADDRD({CLBLM_L_X12Y138_SLICE_X17Y138_BO6, CLBLM_L_X10Y140_SLICE_X12Y140_CO6, CLBLM_R_X11Y138_SLICE_X15Y138_DO6, CLBLM_L_X8Y138_SLICE_X11Y138_DO6, CLBLM_L_X10Y140_SLICE_X13Y140_DO6, CLBLM_R_X11Y139_SLICE_X15Y139_DO6}),
.DIA(CLBLM_L_X10Y139_SLICE_X13Y139_BO6),
.DIB(CLBLM_R_X13Y142_SLICE_X18Y142_AO6),
.DIC(CLBLM_R_X13Y141_SLICE_X18Y141_CO6),
.DID(1'b0),
.DOA(CLBLM_R_X13Y140_SLICE_X18Y140_AO6),
.DOB(CLBLM_R_X13Y140_SLICE_X18Y140_BO6),
.DOC(CLBLM_R_X13Y140_SLICE_X18Y140_CO6),
.DOD(CLBLM_R_X13Y140_SLICE_X18Y140_DO6),
.WCLK(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.WE(CLBLM_L_X12Y139_SLICE_X17Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_DO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_CO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa5555fffff0f0)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_BO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c0000000400000)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLM_R_X13Y138_SLICE_X19Y138_DO6),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_DO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccceccccccc)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_L_X12Y141_SLICE_X17Y141_CO6),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_CO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0040ffff0000)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I4(CLBLM_R_X13Y141_SLICE_X18Y141_AO6),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cf808fc0cfc0cf)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_ALUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_BO6),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.Q(CLBLM_R_X13Y141_SLICE_X19Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_R_X13Y141_SLICE_X19Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_R_X13Y141_SLICE_X19Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_DO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f7f70000d5d5)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_CLUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_BO6),
.I1(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I2(CLBLM_R_X15Y143_SLICE_X20Y143_DO6),
.I3(1'b1),
.I4(CLBLM_R_X15Y139_SLICE_X20Y139_AO6),
.I5(CLBLM_R_X13Y141_SLICE_X19Y141_BO6),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_CO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033550fff33550f)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_BLUT (
.I0(CLBLM_R_X15Y142_SLICE_X21Y142_DQ),
.I1(CLBLM_R_X15Y141_SLICE_X21Y141_BQ),
.I2(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I5(CLBLM_L_X16Y142_SLICE_X22Y142_CQ),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_BO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_AO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_DO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_CO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55f35500550055)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_BLUT (
.I0(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_AO5),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_BO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff08ff00ff00)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_A5Q),
.I3(CLBLM_R_X13Y142_SLICE_X18Y142_BO6),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_AO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_DO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_CO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_BO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_AO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X13Y144_SLICE_X18Y144_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X13Y144_SLICE_X18Y144_D_CY, CLBLM_R_X13Y144_SLICE_X18Y144_C_CY, CLBLM_R_X13Y144_SLICE_X18Y144_B_CY, CLBLM_R_X13Y144_SLICE_X18Y144_A_CY}),
.CYINIT(CLBLM_L_X12Y144_SLICE_X16Y144_DO6),
.DI({1'b0, 1'b0, 1'b0, CLBLM_R_X13Y144_SLICE_X18Y144_AO5}),
.O({CLBLM_R_X13Y144_SLICE_X18Y144_D_XOR, CLBLM_R_X13Y144_SLICE_X18Y144_C_XOR, CLBLM_R_X13Y144_SLICE_X18Y144_B_XOR, CLBLM_R_X13Y144_SLICE_X18Y144_A_XOR}),
.S({CLBLM_R_X13Y144_SLICE_X18Y144_DO6, CLBLM_R_X13Y144_SLICE_X18Y144_CO6, CLBLM_R_X13Y144_SLICE_X18Y144_BO6, CLBLM_R_X13Y144_SLICE_X18Y144_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_DLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_DO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_CO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_BO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00000000)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_AO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00055553333)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_DLUT (
.I0(CLBLM_R_X13Y144_SLICE_X18Y144_D_XOR),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_DO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33553355fff000f0)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_A_XOR),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I4(CLBLM_R_X13Y145_SLICE_X18Y145_B_XOR),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_CO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd3cfd3cec3cec3c)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_BO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77334433440077)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_ALUT (
.I0(CLBLM_R_X13Y145_SLICE_X19Y145_BO5),
.I1(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_AO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X13Y144_SLICE_X19Y144_MUXF7A (
.I0(CLBLM_R_X13Y144_SLICE_X19Y144_BO6),
.I1(CLBLM_R_X13Y144_SLICE_X19Y144_AO6),
.O(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.S(CLBLM_R_X15Y146_SLICE_X20Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X13Y145_SLICE_X18Y145_CARRY4 (
.CI(CLBLM_R_X13Y144_SLICE_X18Y144_COUT),
.CO({CLBLM_R_X13Y145_SLICE_X18Y145_D_CY, CLBLM_R_X13Y145_SLICE_X18Y145_C_CY, CLBLM_R_X13Y145_SLICE_X18Y145_B_CY, CLBLM_R_X13Y145_SLICE_X18Y145_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X13Y145_SLICE_X18Y145_D_XOR, CLBLM_R_X13Y145_SLICE_X18Y145_C_XOR, CLBLM_R_X13Y145_SLICE_X18Y145_B_XOR, CLBLM_R_X13Y145_SLICE_X18Y145_A_XOR}),
.S({CLBLM_R_X13Y145_SLICE_X18Y145_DO6, CLBLM_R_X13Y145_SLICE_X18Y145_CO6, CLBLM_R_X13Y145_SLICE_X18Y145_BO6, CLBLM_R_X13Y145_SLICE_X18Y145_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_DO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_CLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_CO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_BO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_AO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_DO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0ffcc3300)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y146_SLICE_X20Y146_AO6),
.I2(CLBLM_R_X13Y144_SLICE_X19Y144_DO6),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_AO6),
.I4(CLBLM_R_X13Y148_SLICE_X18Y148_AO6),
.I5(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_CO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ee22ee22)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I2(CLBLM_R_X13Y145_SLICE_X18Y145_C_XOR),
.I3(CLBLM_R_X13Y145_SLICE_X18Y145_A_XOR),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_BO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfffb0805f505f5)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I4(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_AO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X13Y146_SLICE_X18Y146_CARRY4 (
.CI(CLBLM_R_X13Y145_SLICE_X18Y145_COUT),
.CO({CLBLM_R_X13Y146_SLICE_X18Y146_D_CY, CLBLM_R_X13Y146_SLICE_X18Y146_C_CY, CLBLM_R_X13Y146_SLICE_X18Y146_B_CY, CLBLM_R_X13Y146_SLICE_X18Y146_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X13Y146_SLICE_X18Y146_D_XOR, CLBLM_R_X13Y146_SLICE_X18Y146_C_XOR, CLBLM_R_X13Y146_SLICE_X18Y146_B_XOR, CLBLM_R_X13Y146_SLICE_X18Y146_A_XOR}),
.S({CLBLM_R_X13Y146_SLICE_X18Y146_DO6, CLBLM_R_X13Y146_SLICE_X18Y146_CO6, CLBLM_R_X13Y146_SLICE_X18Y146_BO6, CLBLM_R_X13Y146_SLICE_X18Y146_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_DO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_CO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_BO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_R_X13Y146_SLICE_X18Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.O5(CLBLM_R_X13Y146_SLICE_X18Y146_AO5),
.O6(CLBLM_R_X13Y146_SLICE_X18Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf88df8888dd88df)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_DO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30500050f050c050)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_CO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000feaabaaa)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_BLUT (
.I0(CLBLM_R_X13Y146_SLICE_X19Y146_DO6),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I5(CLBLM_R_X13Y146_SLICE_X19Y146_CO6),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_BO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4200440000001000)
  ) CLBLM_R_X13Y146_SLICE_X19Y146_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y146_SLICE_X19Y146_AO5),
.O6(CLBLM_R_X13Y146_SLICE_X19Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X13Y147_SLICE_X18Y147_CARRY4 (
.CI(CLBLM_R_X13Y146_SLICE_X18Y146_COUT),
.CO({CLBLM_R_X13Y147_SLICE_X18Y147_D_CY, CLBLM_R_X13Y147_SLICE_X18Y147_C_CY, CLBLM_R_X13Y147_SLICE_X18Y147_B_CY, CLBLM_R_X13Y147_SLICE_X18Y147_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X13Y147_SLICE_X18Y147_D_XOR, CLBLM_R_X13Y147_SLICE_X18Y147_C_XOR, CLBLM_R_X13Y147_SLICE_X18Y147_B_XOR, CLBLM_R_X13Y147_SLICE_X18Y147_A_XOR}),
.S({CLBLM_R_X13Y147_SLICE_X18Y147_DO6, CLBLM_R_X13Y147_SLICE_X18Y147_CO6, CLBLM_R_X13Y147_SLICE_X18Y147_BO6, CLBLM_R_X13Y147_SLICE_X18Y147_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_DO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_CO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_BO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_AO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heecceccccccceccc)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_R_X13Y146_SLICE_X19Y146_DO6),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_DO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1104110411550044)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_CLUT (
.I0(CLBLM_R_X13Y147_SLICE_X19Y147_AO6),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I4(CLBLM_L_X16Y152_SLICE_X23Y152_AO6),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_CO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff08ccffff19dd)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_BLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I2(CLBLM_R_X13Y148_SLICE_X19Y148_DO6),
.I3(CLBLM_R_X13Y147_SLICE_X19Y147_DO6),
.I4(CLBLM_R_X13Y147_SLICE_X19Y147_CO6),
.I5(CLBLM_R_X13Y148_SLICE_X19Y148_CO6),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_BO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ffff0005ffff)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_DLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_BO5),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_DO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a0003333b333)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I4(CLBLM_R_X13Y148_SLICE_X18Y148_DO6),
.I5(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_CO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacc0cf00000000)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_BLUT (
.I0(CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR),
.I1(CLBLM_R_X15Y148_SLICE_X21Y148_AO6),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_BO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcccc3366669999)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_AO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7807700ff887f08)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_DO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cec16b616b64cec)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_CLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I3(CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_CO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffdff00ffff)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_BLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I1(CLBLM_R_X13Y149_SLICE_X19Y149_AO6),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I4(CLBLM_R_X13Y148_SLICE_X19Y148_AO6),
.I5(CLBLM_R_X13Y149_SLICE_X19Y149_AO5),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_BO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1020ffffffffffff)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_AO6),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_AO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffcc)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR),
.I2(1'b1),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_DO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9633333396333333)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_CLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_CO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddf5ffff88a00000)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR),
.I2(CLBLM_R_X13Y148_SLICE_X18Y148_AO5),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_R_X13Y149_SLICE_X18Y149_CO6),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_BO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f2c2f2c1310d3d0)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_ALUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I3(CLBLM_R_X15Y153_SLICE_X21Y153_CO6),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_AO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X13Y149_SLICE_X18Y149_MUXF7A (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_BO6),
.I1(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.O(CLBLM_R_X13Y149_SLICE_X18Y149_F7AMUX_O),
.S(CLBLM_R_X15Y150_SLICE_X20Y150_DO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_DO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_CO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_BO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44404040bbbebebe)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_ALUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_AO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5353535353535353)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_DO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f7766660f666666)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_CO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bcf0f0f8b030f0f)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_BLUT (
.I0(CLBLM_R_X13Y150_SLICE_X18Y150_DO6),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_R_X13Y144_SLICE_X19Y144_CO5),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_BO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50eeeefa504444)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_ALUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_BO6),
.I2(CLBLM_R_X15Y150_SLICE_X21Y150_BO6),
.I3(CLBLM_R_X13Y150_SLICE_X18Y150_BO6),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I5(CLBLM_R_X13Y150_SLICE_X18Y150_CO6),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_AO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505955505056555)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_DLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_DO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ccc5dffa200a200)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_CO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaaeaaabaaaaaaa)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_BLUT (
.I0(CLBLM_R_X13Y150_SLICE_X19Y150_DO6),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.I5(CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_BO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5757f5a00202f5a0)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I3(CLBLM_R_X15Y151_SLICE_X20Y151_CO5),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(CLBLM_R_X13Y150_SLICE_X19Y150_CO6),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_AO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X13Y150_SLICE_X19Y150_MUXF7A (
.I0(CLBLM_R_X13Y150_SLICE_X19Y150_BO6),
.I1(CLBLM_R_X13Y150_SLICE_X19Y150_AO6),
.O(CLBLM_R_X13Y150_SLICE_X19Y150_F7AMUX_O),
.S(CLBLM_R_X15Y150_SLICE_X20Y150_DO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y128_SLICE_X20Y128_AO5),
.Q(CLBLM_R_X15Y128_SLICE_X20Y128_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y128_SLICE_X20Y128_BO5),
.Q(CLBLM_R_X15Y128_SLICE_X20Y128_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y128_SLICE_X20Y128_AO6),
.Q(CLBLM_R_X15Y128_SLICE_X20Y128_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y128_SLICE_X20Y128_BO6),
.Q(CLBLM_R_X15Y128_SLICE_X20Y128_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y128_SLICE_X20Y128_CO6),
.Q(CLBLM_R_X15Y128_SLICE_X20Y128_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_DO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333333)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_CO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1c1ccccc4a4aaaaa)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_BLUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_B5Q),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_BQ),
.I2(CLBLM_R_X15Y128_SLICE_X20Y128_CQ),
.I3(1'b1),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_BO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200000000ffff00)
  ) CLBLM_R_X15Y128_SLICE_X20Y128_ALUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_B5Q),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_BQ),
.I2(1'b1),
.I3(CLBLM_R_X15Y128_SLICE_X20Y128_CQ),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X20Y128_AO5),
.O6(CLBLM_R_X15Y128_SLICE_X20Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_DO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_CO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_BO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y128_SLICE_X21Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y128_SLICE_X21Y128_AO5),
.O6(CLBLM_R_X15Y128_SLICE_X21Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y129_SLICE_X20Y129_AO6),
.Q(CLBLM_R_X15Y129_SLICE_X20Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y129_SLICE_X20Y129_BO6),
.Q(CLBLM_R_X15Y129_SLICE_X20Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y129_SLICE_X20Y129_CO6),
.Q(CLBLM_R_X15Y129_SLICE_X20Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_DO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafffafffafffbfbf)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_CLUT (
.I0(CLBLM_R_X15Y131_SLICE_X20Y131_AQ),
.I1(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I2(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_CO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f7fffdffff)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_BLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLM_R_X15Y129_SLICE_X20Y129_CQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_BO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddffffdffff)
  ) CLBLM_R_X15Y129_SLICE_X20Y129_ALUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I1(CLBLM_R_X15Y129_SLICE_X20Y129_BQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.O5(CLBLM_R_X15Y129_SLICE_X20Y129_AO5),
.O6(CLBLM_R_X15Y129_SLICE_X20Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y129_SLICE_X21Y129_BO5),
.Q(CLBLM_R_X15Y129_SLICE_X21Y129_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y129_SLICE_X21Y129_AO6),
.Q(CLBLM_R_X15Y129_SLICE_X21Y129_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y129_SLICE_X21Y129_BO6),
.Q(CLBLM_R_X15Y129_SLICE_X21Y129_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y129_SLICE_X21Y129_CO6),
.Q(CLBLM_R_X15Y129_SLICE_X21Y129_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003000000030)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y129_SLICE_X21Y129_CQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_DO6),
.I3(CLBLM_R_X15Y130_SLICE_X21Y130_DO6),
.I4(CLBLM_R_X15Y129_SLICE_X21Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_DO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff05f5cccccccc)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_CLUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I1(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I3(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_CO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f044f0ff000000)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_BLUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I2(CLBLM_R_X15Y129_SLICE_X21Y129_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_BO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30b830fc30fc74)
  ) CLBLM_R_X15Y129_SLICE_X21Y129_ALUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I2(CLBLM_R_X15Y129_SLICE_X21Y129_CQ),
.I3(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.O5(CLBLM_R_X15Y129_SLICE_X21Y129_AO5),
.O6(CLBLM_R_X15Y129_SLICE_X21Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y130_SLICE_X20Y130_AO6),
.D(LIOB33_X0Y101_IOB_X0Y101_I),
.PRE(LIOB33_X0Y105_IOB_X0Y106_I),
.Q(CLBLM_R_X15Y130_SLICE_X20Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_DO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_CO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_BO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000050500000303)
  ) CLBLM_R_X15Y130_SLICE_X20Y130_ALUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I1(CLBLM_R_X13Y136_SLICE_X19Y136_BQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_BO6),
.I3(1'b1),
.I4(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.O5(CLBLM_R_X15Y130_SLICE_X20Y130_AO5),
.O6(CLBLM_R_X15Y130_SLICE_X20Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y130_SLICE_X21Y130_AO6),
.Q(CLBLM_R_X15Y130_SLICE_X21Y130_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y130_SLICE_X21Y130_BO6),
.Q(CLBLM_R_X15Y130_SLICE_X21Y130_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y130_SLICE_X21Y130_CO6),
.Q(CLBLM_R_X15Y130_SLICE_X21Y130_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffc)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y130_SLICE_X21Y130_CQ),
.I2(CLBLM_L_X16Y131_SLICE_X22Y131_AQ),
.I3(CLBLM_R_X15Y130_SLICE_X21Y130_BQ),
.I4(CLBLM_R_X15Y130_SLICE_X21Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_DO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555533f0f0f0f0)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_CLUT (
.I0(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I1(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I2(CLBLM_L_X16Y131_SLICE_X22Y131_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_CO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f033f022f077f0)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_BLUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I1(CLBLM_R_X15Y144_SLICE_X21Y144_CO6),
.I2(CLBLM_R_X15Y130_SLICE_X21Y130_CQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I4(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_BO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05ccffcc00ccfacc)
  ) CLBLM_R_X15Y130_SLICE_X21Y130_ALUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I1(CLBLM_R_X15Y130_SLICE_X21Y130_BQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.O5(CLBLM_R_X15Y130_SLICE_X21Y130_AO5),
.O6(CLBLM_R_X15Y130_SLICE_X21Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y131_SLICE_X20Y131_AO6),
.Q(CLBLM_R_X15Y131_SLICE_X20Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y131_SLICE_X20Y131_BO6),
.Q(CLBLM_R_X15Y131_SLICE_X20Y131_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y131_SLICE_X20Y131_CO6),
.Q(CLBLM_R_X15Y131_SLICE_X20Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y130_SLICE_X18Y130_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y131_SLICE_X20Y131_DO6),
.Q(CLBLM_R_X15Y131_SLICE_X20Y131_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff01fdffff)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_DLUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I5(CLBLM_R_X13Y131_SLICE_X19Y131_BQ),
.O5(CLBLM_R_X15Y131_SLICE_X20Y131_DO5),
.O6(CLBLM_R_X15Y131_SLICE_X20Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fffffff1fdffff)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_CLUT (
.I0(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_DQ),
.I3(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.I4(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.O5(CLBLM_R_X15Y131_SLICE_X20Y131_CO5),
.O6(CLBLM_R_X15Y131_SLICE_X20Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f7fffdffff)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_BLUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_CQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.O5(CLBLM_R_X15Y131_SLICE_X20Y131_BO5),
.O6(CLBLM_R_X15Y131_SLICE_X20Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddffffdffff)
  ) CLBLM_R_X15Y131_SLICE_X20Y131_ALUT (
.I0(CLBLM_R_X13Y130_SLICE_X19Y130_AQ),
.I1(CLBLM_R_X15Y131_SLICE_X20Y131_BQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I4(CLBLM_R_X15Y128_SLICE_X20Y128_AQ),
.I5(CLBLM_R_X13Y132_SLICE_X18Y132_DQ),
.O5(CLBLM_R_X15Y131_SLICE_X20Y131_AO5),
.O6(CLBLM_R_X15Y131_SLICE_X20Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y131_SLICE_X21Y131_BO5),
.Q(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y131_SLICE_X21Y131_AO6),
.Q(CLBLM_R_X15Y131_SLICE_X21Y131_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X12Y129_SLICE_X17Y129_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y131_SLICE_X21Y131_CO6),
.Q(CLBLM_R_X15Y131_SLICE_X21Y131_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000003)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y131_SLICE_X21Y131_CQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I3(CLBLM_R_X15Y129_SLICE_X21Y129_B5Q),
.I4(CLBLM_R_X15Y131_SLICE_X21Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y131_SLICE_X21Y131_DO5),
.O6(CLBLM_R_X15Y131_SLICE_X21Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0a5f0a5f0a7722)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I3(CLBLM_R_X15Y131_SLICE_X21Y131_A5Q),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.O5(CLBLM_R_X15Y131_SLICE_X21Y131_CO5),
.O6(CLBLM_R_X15Y131_SLICE_X21Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h003300335577f0f0)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_BLUT (
.I0(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I2(CLBLM_R_X15Y131_SLICE_X21Y131_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y131_SLICE_X21Y131_BO5),
.O6(CLBLM_R_X15Y131_SLICE_X21Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acacacaca)
  ) CLBLM_R_X15Y131_SLICE_X21Y131_ALUT (
.I0(CLBLM_R_X15Y129_SLICE_X21Y129_B5Q),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BQ),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I3(1'b1),
.I4(CLBLM_R_X13Y136_SLICE_X19Y136_AQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.O5(CLBLM_R_X15Y131_SLICE_X21Y131_AO5),
.O6(CLBLM_R_X15Y131_SLICE_X21Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y133_SLICE_X20Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y133_SLICE_X20Y133_DO5),
.O6(CLBLM_R_X15Y133_SLICE_X20Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y133_SLICE_X20Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y133_SLICE_X20Y133_CO5),
.O6(CLBLM_R_X15Y133_SLICE_X20Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y133_SLICE_X20Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y133_SLICE_X20Y133_BO5),
.O6(CLBLM_R_X15Y133_SLICE_X20Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y133_SLICE_X20Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y133_SLICE_X20Y133_AO5),
.O6(CLBLM_R_X15Y133_SLICE_X20Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y133_SLICE_X21Y133_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y133_SLICE_X21Y133_AO6),
.Q(CLBLM_R_X15Y133_SLICE_X21Y133_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y133_SLICE_X21Y133_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y133_SLICE_X21Y133_BO6),
.Q(CLBLM_R_X15Y133_SLICE_X21Y133_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y133_SLICE_X21Y133_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y133_SLICE_X21Y133_CO6),
.Q(CLBLM_R_X15Y133_SLICE_X21Y133_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y133_SLICE_X21Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y133_SLICE_X21Y133_DO5),
.O6(CLBLM_R_X15Y133_SLICE_X21Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030fcfc2230eefc)
  ) CLBLM_R_X15Y133_SLICE_X21Y133_CLUT (
.I0(CLBLM_R_X15Y134_SLICE_X20Y134_D_XOR),
.I1(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.I2(CLBLM_R_X13Y133_SLICE_X19Y133_B5Q),
.I3(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I4(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O5(CLBLM_R_X15Y133_SLICE_X21Y133_CO5),
.O6(CLBLM_R_X15Y133_SLICE_X21Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcc0faa0fcc0fcc)
  ) CLBLM_R_X15Y133_SLICE_X21Y133_BLUT (
.I0(CLBLM_R_X15Y134_SLICE_X20Y134_B_XOR),
.I1(CLBLM_R_X13Y133_SLICE_X19Y133_BQ),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I3(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I5(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.O5(CLBLM_R_X15Y133_SLICE_X21Y133_BO5),
.O6(CLBLM_R_X15Y133_SLICE_X21Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf055ccccf0f0)
  ) CLBLM_R_X15Y133_SLICE_X21Y133_ALUT (
.I0(CLBLM_R_X15Y133_SLICE_X21Y133_AQ),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I2(CLBLM_R_X13Y133_SLICE_X19Y133_AQ),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I4(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.I5(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.O5(CLBLM_R_X15Y133_SLICE_X21Y133_AO5),
.O6(CLBLM_R_X15Y133_SLICE_X21Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y134_SLICE_X20Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y134_SLICE_X20Y134_BO5),
.Q(CLBLM_R_X15Y134_SLICE_X20Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y134_SLICE_X20Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y134_SLICE_X20Y134_CO5),
.Q(CLBLM_R_X15Y134_SLICE_X20Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y134_SLICE_X20Y134_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y129_SLICE_X19Y129_AQ),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y134_SLICE_X20Y134_DO5),
.Q(CLBLM_R_X15Y134_SLICE_X20Y134_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X15Y134_SLICE_X20Y134_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X15Y134_SLICE_X20Y134_D_CY, CLBLM_R_X15Y134_SLICE_X20Y134_C_CY, CLBLM_R_X15Y134_SLICE_X20Y134_B_CY, CLBLM_R_X15Y134_SLICE_X20Y134_A_CY}),
.CYINIT(CLBLM_R_X15Y133_SLICE_X21Y133_AQ),
.DI({1'b0, 1'b0, 1'b0, CLBLM_R_X15Y134_SLICE_X20Y134_AO5}),
.O({CLBLM_R_X15Y134_SLICE_X20Y134_D_XOR, CLBLM_R_X15Y134_SLICE_X20Y134_C_XOR, CLBLM_R_X15Y134_SLICE_X20Y134_B_XOR, CLBLM_R_X15Y134_SLICE_X20Y134_A_XOR}),
.S({CLBLM_R_X15Y134_SLICE_X20Y134_DO6, CLBLM_R_X15Y134_SLICE_X20Y134_CO6, CLBLM_R_X15Y134_SLICE_X20Y134_BO6, CLBLM_R_X15Y134_SLICE_X20Y134_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00ff00)
  ) CLBLM_R_X15Y134_SLICE_X20Y134_DLUT (
.I0(CLBLM_R_X15Y133_SLICE_X21Y133_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y134_SLICE_X20Y134_DO5),
.O6(CLBLM_R_X15Y134_SLICE_X20Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_R_X15Y134_SLICE_X20Y134_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y134_SLICE_X21Y134_BQ),
.I2(1'b1),
.I3(CLBLM_R_X15Y131_SLICE_X20Y131_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y134_SLICE_X20Y134_CO5),
.O6(CLBLM_R_X15Y134_SLICE_X20Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0f0f0f0)
  ) CLBLM_R_X15Y134_SLICE_X20Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X15Y131_SLICE_X20Y131_BQ),
.I3(1'b1),
.I4(CLBLM_R_X15Y133_SLICE_X21Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y134_SLICE_X20Y134_BO5),
.O6(CLBLM_R_X15Y134_SLICE_X20Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLM_R_X15Y134_SLICE_X20Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X15Y134_SLICE_X21Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y134_SLICE_X20Y134_AO5),
.O6(CLBLM_R_X15Y134_SLICE_X20Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y134_SLICE_X21Y134_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y134_SLICE_X21Y134_AO6),
.Q(CLBLM_R_X15Y134_SLICE_X21Y134_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y134_SLICE_X21Y134_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y134_SLICE_X21Y134_BO6),
.Q(CLBLM_R_X15Y134_SLICE_X21Y134_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y134_SLICE_X21Y134_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y134_SLICE_X21Y134_CO6),
.Q(CLBLM_R_X15Y134_SLICE_X21Y134_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ffffff77ffffff)
  ) CLBLM_R_X15Y134_SLICE_X21Y134_DLUT (
.I0(CLBLM_R_X15Y135_SLICE_X21Y135_AQ),
.I1(CLBLM_R_X15Y136_SLICE_X21Y136_CQ),
.I2(1'b1),
.I3(CLBLM_R_X15Y134_SLICE_X21Y134_BQ),
.I4(CLBLM_R_X15Y134_SLICE_X21Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y134_SLICE_X21Y134_DO5),
.O6(CLBLM_R_X15Y134_SLICE_X21Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777774744447444)
  ) CLBLM_R_X15Y134_SLICE_X21Y134_CLUT (
.I0(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I1(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.I2(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I3(CLBLM_R_X15Y135_SLICE_X20Y135_A_XOR),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I5(CLBLM_R_X13Y134_SLICE_X19Y134_BQ),
.O5(CLBLM_R_X15Y134_SLICE_X21Y134_CO5),
.O6(CLBLM_R_X15Y134_SLICE_X21Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdff2000fd0020)
  ) CLBLM_R_X15Y134_SLICE_X21Y134_BLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I1(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I2(CLBLM_R_X15Y134_SLICE_X20Y134_C_XOR),
.I3(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.I4(CLBLM_R_X13Y133_SLICE_X19Y133_A5Q),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.O5(CLBLM_R_X15Y134_SLICE_X21Y134_BO5),
.O6(CLBLM_R_X15Y134_SLICE_X21Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fb0008fffbff08)
  ) CLBLM_R_X15Y134_SLICE_X21Y134_ALUT (
.I0(CLBLM_R_X15Y134_SLICE_X20Y134_A_XOR),
.I1(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I2(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I3(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.I4(CLBLM_R_X13Y134_SLICE_X19Y134_AQ),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.O5(CLBLM_R_X15Y134_SLICE_X21Y134_AO5),
.O6(CLBLM_R_X15Y134_SLICE_X21Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X15Y135_SLICE_X20Y135_CARRY4 (
.CI(CLBLM_R_X15Y134_SLICE_X20Y134_COUT),
.CO({CLBLM_R_X15Y135_SLICE_X20Y135_D_CY, CLBLM_R_X15Y135_SLICE_X20Y135_C_CY, CLBLM_R_X15Y135_SLICE_X20Y135_B_CY, CLBLM_R_X15Y135_SLICE_X20Y135_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X15Y135_SLICE_X20Y135_D_XOR, CLBLM_R_X15Y135_SLICE_X20Y135_C_XOR, CLBLM_R_X15Y135_SLICE_X20Y135_B_XOR, CLBLM_R_X15Y135_SLICE_X20Y135_A_XOR}),
.S({CLBLM_R_X15Y135_SLICE_X20Y135_DO6, CLBLM_R_X15Y135_SLICE_X20Y135_CO6, CLBLM_R_X15Y135_SLICE_X20Y135_BO6, CLBLM_R_X15Y135_SLICE_X20Y135_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y135_SLICE_X20Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y136_SLICE_X21Y136_AQ),
.O5(CLBLM_R_X15Y135_SLICE_X20Y135_DO5),
.O6(CLBLM_R_X15Y135_SLICE_X20Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y135_SLICE_X20Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y135_SLICE_X21Y135_BQ),
.O5(CLBLM_R_X15Y135_SLICE_X20Y135_CO5),
.O6(CLBLM_R_X15Y135_SLICE_X20Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y135_SLICE_X20Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y135_SLICE_X21Y135_AQ),
.O5(CLBLM_R_X15Y135_SLICE_X20Y135_BO5),
.O6(CLBLM_R_X15Y135_SLICE_X20Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y135_SLICE_X20Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y134_SLICE_X21Y134_CQ),
.O5(CLBLM_R_X15Y135_SLICE_X20Y135_AO5),
.O6(CLBLM_R_X15Y135_SLICE_X20Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y135_SLICE_X21Y135_AO6),
.Q(CLBLM_R_X15Y135_SLICE_X21Y135_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y135_SLICE_X21Y135_BO6),
.Q(CLBLM_R_X15Y135_SLICE_X21Y135_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccffaaffaa)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_DLUT (
.I0(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.I1(CLBLM_R_X13Y133_SLICE_X19Y133_CO6),
.I2(1'b1),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y135_SLICE_X21Y135_DO5),
.O6(CLBLM_R_X15Y135_SLICE_X21Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdfffffffffffff)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_CLUT (
.I0(CLBLM_R_X15Y136_SLICE_X21Y136_AQ),
.I1(CLBLM_R_X15Y134_SLICE_X21Y134_DO6),
.I2(CLBLM_R_X15Y138_SLICE_X21Y138_BQ),
.I3(1'b1),
.I4(CLBLM_R_X15Y136_SLICE_X21Y136_DQ),
.I5(CLBLM_R_X15Y137_SLICE_X21Y137_BQ),
.O5(CLBLM_R_X15Y135_SLICE_X21Y135_CO5),
.O6(CLBLM_R_X15Y135_SLICE_X21Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fd20fffffd20)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_BLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I1(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I2(CLBLM_R_X15Y135_SLICE_X20Y135_C_XOR),
.I3(CLBLM_R_X13Y134_SLICE_X19Y134_A5Q),
.I4(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.I5(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.O5(CLBLM_R_X15Y135_SLICE_X21Y135_BO5),
.O6(CLBLM_R_X15Y135_SLICE_X21Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0e0c04fcfefcf4)
  ) CLBLM_R_X15Y135_SLICE_X21Y135_ALUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I1(CLBLM_R_X13Y134_SLICE_X19Y134_B5Q),
.I2(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I4(CLBLM_R_X15Y135_SLICE_X20Y135_B_XOR),
.I5(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.O5(CLBLM_R_X15Y135_SLICE_X21Y135_AO5),
.O6(CLBLM_R_X15Y135_SLICE_X21Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X15Y136_SLICE_X20Y136_CARRY4 (
.CI(CLBLM_R_X15Y135_SLICE_X20Y135_COUT),
.CO({CLBLM_R_X15Y136_SLICE_X20Y136_D_CY, CLBLM_R_X15Y136_SLICE_X20Y136_C_CY, CLBLM_R_X15Y136_SLICE_X20Y136_B_CY, CLBLM_R_X15Y136_SLICE_X20Y136_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X15Y136_SLICE_X20Y136_D_XOR, CLBLM_R_X15Y136_SLICE_X20Y136_C_XOR, CLBLM_R_X15Y136_SLICE_X20Y136_B_XOR, CLBLM_R_X15Y136_SLICE_X20Y136_A_XOR}),
.S({CLBLM_R_X15Y136_SLICE_X20Y136_DO6, CLBLM_R_X15Y136_SLICE_X20Y136_CO6, CLBLM_R_X15Y136_SLICE_X20Y136_BO6, CLBLM_R_X15Y136_SLICE_X20Y136_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y136_SLICE_X20Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y136_SLICE_X21Y136_DQ),
.O5(CLBLM_R_X15Y136_SLICE_X20Y136_DO5),
.O6(CLBLM_R_X15Y136_SLICE_X20Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y136_SLICE_X20Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y136_SLICE_X21Y136_CQ),
.O5(CLBLM_R_X15Y136_SLICE_X20Y136_CO5),
.O6(CLBLM_R_X15Y136_SLICE_X20Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y136_SLICE_X20Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y136_SLICE_X21Y136_BQ),
.O5(CLBLM_R_X15Y136_SLICE_X20Y136_BO5),
.O6(CLBLM_R_X15Y136_SLICE_X20Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y136_SLICE_X20Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y137_SLICE_X21Y137_AQ),
.O5(CLBLM_R_X15Y136_SLICE_X20Y136_AO5),
.O6(CLBLM_R_X15Y136_SLICE_X20Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y136_SLICE_X21Y136_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y136_SLICE_X21Y136_AO6),
.Q(CLBLM_R_X15Y136_SLICE_X21Y136_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y136_SLICE_X21Y136_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y136_SLICE_X21Y136_BO6),
.Q(CLBLM_R_X15Y136_SLICE_X21Y136_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y136_SLICE_X21Y136_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y136_SLICE_X21Y136_CO6),
.Q(CLBLM_R_X15Y136_SLICE_X21Y136_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y136_SLICE_X21Y136_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y136_SLICE_X21Y136_DO6),
.Q(CLBLM_R_X15Y136_SLICE_X21Y136_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffba8aba8a)
  ) CLBLM_R_X15Y136_SLICE_X21Y136_DLUT (
.I0(CLBLM_R_X13Y136_SLICE_X18Y136_B5Q),
.I1(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I2(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I3(CLBLM_R_X15Y136_SLICE_X20Y136_D_XOR),
.I4(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I5(CLBLM_R_X13Y133_SLICE_X19Y133_CO6),
.O5(CLBLM_R_X15Y136_SLICE_X21Y136_DO5),
.O6(CLBLM_R_X15Y136_SLICE_X21Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5e4e4e4a0e4e4)
  ) CLBLM_R_X15Y136_SLICE_X21Y136_CLUT (
.I0(CLBLM_R_X13Y133_SLICE_X19Y133_CO6),
.I1(CLBLM_R_X13Y136_SLICE_X18Y136_A5Q),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I4(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I5(CLBLM_R_X15Y136_SLICE_X20Y136_C_XOR),
.O5(CLBLM_R_X15Y136_SLICE_X21Y136_CO5),
.O6(CLBLM_R_X15Y136_SLICE_X21Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fcccc0f0fee44)
  ) CLBLM_R_X15Y136_SLICE_X21Y136_BLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I1(CLBLM_R_X13Y136_SLICE_X18Y136_BQ),
.I2(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I3(CLBLM_R_X15Y136_SLICE_X20Y136_B_XOR),
.I4(CLBLM_R_X13Y133_SLICE_X19Y133_CO6),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O5(CLBLM_R_X15Y136_SLICE_X21Y136_BO5),
.O6(CLBLM_R_X15Y136_SLICE_X21Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffddf0f02200)
  ) CLBLM_R_X15Y136_SLICE_X21Y136_ALUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I1(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I3(CLBLM_R_X15Y135_SLICE_X20Y135_D_XOR),
.I4(CLBLM_R_X13Y133_SLICE_X19Y133_CO6),
.I5(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.O5(CLBLM_R_X15Y136_SLICE_X21Y136_AO5),
.O6(CLBLM_R_X15Y136_SLICE_X21Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X15Y137_SLICE_X20Y137_CARRY4 (
.CI(CLBLM_R_X15Y136_SLICE_X20Y136_COUT),
.CO({CLBLM_R_X15Y137_SLICE_X20Y137_D_CY, CLBLM_R_X15Y137_SLICE_X20Y137_C_CY, CLBLM_R_X15Y137_SLICE_X20Y137_B_CY, CLBLM_R_X15Y137_SLICE_X20Y137_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X15Y137_SLICE_X20Y137_D_XOR, CLBLM_R_X15Y137_SLICE_X20Y137_C_XOR, CLBLM_R_X15Y137_SLICE_X20Y137_B_XOR, CLBLM_R_X15Y137_SLICE_X20Y137_A_XOR}),
.S({CLBLM_R_X15Y137_SLICE_X20Y137_DO6, CLBLM_R_X15Y137_SLICE_X20Y137_CO6, CLBLM_R_X15Y137_SLICE_X20Y137_BO6, CLBLM_R_X15Y137_SLICE_X20Y137_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffff)
  ) CLBLM_R_X15Y137_SLICE_X20Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y137_SLICE_X20Y137_DO5),
.O6(CLBLM_R_X15Y137_SLICE_X20Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y137_SLICE_X20Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y138_SLICE_X21Y138_BQ),
.O5(CLBLM_R_X15Y137_SLICE_X20Y137_CO5),
.O6(CLBLM_R_X15Y137_SLICE_X20Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y137_SLICE_X20Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y138_SLICE_X21Y138_AQ),
.O5(CLBLM_R_X15Y137_SLICE_X20Y137_BO5),
.O6(CLBLM_R_X15Y137_SLICE_X20Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y137_SLICE_X20Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y137_SLICE_X21Y137_BQ),
.O5(CLBLM_R_X15Y137_SLICE_X20Y137_AO5),
.O6(CLBLM_R_X15Y137_SLICE_X20Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y137_SLICE_X21Y137_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y137_SLICE_X21Y137_AO6),
.Q(CLBLM_R_X15Y137_SLICE_X21Y137_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y137_SLICE_X21Y137_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y137_SLICE_X21Y137_BO6),
.Q(CLBLM_R_X15Y137_SLICE_X21Y137_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h04340737c4f4c7f7)
  ) CLBLM_R_X15Y137_SLICE_X21Y137_DLUT (
.I0(CLBLM_R_X15Y134_SLICE_X20Y134_CQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.I3(CLBLM_L_X16Y136_SLICE_X23Y136_AQ),
.I4(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I5(CLBLL_L_X26Y135_SLICE_X38Y135_AO6),
.O5(CLBLM_R_X15Y137_SLICE_X21Y137_DO5),
.O6(CLBLM_R_X15Y137_SLICE_X21Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeeefe00044404)
  ) CLBLM_R_X15Y137_SLICE_X21Y137_CLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.I1(CLBLL_L_X26Y135_SLICE_X38Y135_AO5),
.I2(CLBLM_R_X15Y142_SLICE_X20Y142_DO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLL_L_X26Y135_SLICE_X38Y135_AO6),
.O5(CLBLM_R_X15Y137_SLICE_X21Y137_CO5),
.O6(CLBLM_R_X15Y137_SLICE_X21Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2e2e2e2e3f0c2e2e)
  ) CLBLM_R_X15Y137_SLICE_X21Y137_BLUT (
.I0(CLBLM_L_X12Y138_SLICE_X17Y138_AQ),
.I1(CLBLM_R_X13Y133_SLICE_X19Y133_CO6),
.I2(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I3(CLBLM_R_X15Y137_SLICE_X20Y137_A_XOR),
.I4(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O5(CLBLM_R_X15Y137_SLICE_X21Y137_BO5),
.O6(CLBLM_R_X15Y137_SLICE_X21Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0c3f0c3f2e1d0c)
  ) CLBLM_R_X15Y137_SLICE_X21Y137_ALUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I1(CLBLM_R_X13Y133_SLICE_X19Y133_CO6),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I3(CLBLM_R_X13Y138_SLICE_X18Y138_AQ),
.I4(CLBLM_R_X15Y136_SLICE_X20Y136_A_XOR),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O5(CLBLM_R_X15Y137_SLICE_X21Y137_AO5),
.O6(CLBLM_R_X15Y137_SLICE_X21Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y138_SLICE_X20Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y138_SLICE_X20Y138_DO5),
.O6(CLBLM_R_X15Y138_SLICE_X20Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y138_SLICE_X20Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y138_SLICE_X20Y138_CO5),
.O6(CLBLM_R_X15Y138_SLICE_X20Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y138_SLICE_X20Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y138_SLICE_X20Y138_BO5),
.O6(CLBLM_R_X15Y138_SLICE_X20Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y138_SLICE_X20Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y138_SLICE_X20Y138_AO5),
.O6(CLBLM_R_X15Y138_SLICE_X20Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y138_SLICE_X21Y138_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y138_SLICE_X21Y138_AO6),
.Q(CLBLM_R_X15Y138_SLICE_X21Y138_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y138_SLICE_X21Y138_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y135_SLICE_X21Y135_DO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y138_SLICE_X21Y138_BO6),
.Q(CLBLM_R_X15Y138_SLICE_X21Y138_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y138_SLICE_X21Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y138_SLICE_X21Y138_DO5),
.O6(CLBLM_R_X15Y138_SLICE_X21Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y138_SLICE_X21Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y138_SLICE_X21Y138_CO5),
.O6(CLBLM_R_X15Y138_SLICE_X21Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f35303a3030)
  ) CLBLM_R_X15Y138_SLICE_X21Y138_BLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I2(CLBLM_R_X13Y133_SLICE_X19Y133_CO6),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I4(CLBLM_R_X15Y137_SLICE_X20Y137_C_XOR),
.I5(CLBLM_R_X13Y138_SLICE_X18Y138_A5Q),
.O5(CLBLM_R_X15Y138_SLICE_X21Y138_BO5),
.O6(CLBLM_R_X15Y138_SLICE_X21Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0d0008fffdf0f8)
  ) CLBLM_R_X15Y138_SLICE_X21Y138_ALUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.I1(CLBLM_R_X15Y137_SLICE_X20Y137_B_XOR),
.I2(CLBLM_R_X13Y133_SLICE_X19Y133_CO6),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I4(CLBLM_L_X12Y138_SLICE_X17Y138_BQ),
.I5(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.O5(CLBLM_R_X15Y138_SLICE_X21Y138_AO5),
.O6(CLBLM_R_X15Y138_SLICE_X21Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y139_SLICE_X20Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y139_SLICE_X20Y139_DO5),
.O6(CLBLM_R_X15Y139_SLICE_X20Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y139_SLICE_X20Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y139_SLICE_X20Y139_CO5),
.O6(CLBLM_R_X15Y139_SLICE_X20Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y139_SLICE_X20Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y139_SLICE_X20Y139_BO5),
.O6(CLBLM_R_X15Y139_SLICE_X20Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000410082)
  ) CLBLM_R_X15Y139_SLICE_X20Y139_ALUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I2(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I3(CLBLM_L_X10Y138_SLICE_X13Y138_BO6),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_CO6),
.O5(CLBLM_R_X15Y139_SLICE_X20Y139_AO5),
.O6(CLBLM_R_X15Y139_SLICE_X20Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y139_SLICE_X21Y139_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_R_X15Y139_SLICE_X21Y139_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y139_SLICE_X21Y139_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_R_X15Y139_SLICE_X21Y139_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y139_SLICE_X21Y139_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_R_X15Y139_SLICE_X21Y139_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y139_SLICE_X21Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y139_SLICE_X21Y139_DO5),
.O6(CLBLM_R_X15Y139_SLICE_X21Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y139_SLICE_X21Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y139_SLICE_X21Y139_CO5),
.O6(CLBLM_R_X15Y139_SLICE_X21Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h11bb0a0a11bb5f5f)
  ) CLBLM_R_X15Y139_SLICE_X21Y139_BLUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I1(CLBLM_L_X16Y140_SLICE_X22Y140_CQ),
.I2(CLBLM_R_X15Y140_SLICE_X21Y140_DQ),
.I3(CLBLM_R_X15Y139_SLICE_X21Y139_CQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(CLBLM_R_X15Y140_SLICE_X20Y140_CQ),
.O5(CLBLM_R_X15Y139_SLICE_X21Y139_BO5),
.O6(CLBLM_R_X15Y139_SLICE_X21Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f440f770f)
  ) CLBLM_R_X15Y139_SLICE_X21Y139_ALUT (
.I0(CLBLM_R_X15Y139_SLICE_X21Y139_BO6),
.I1(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I2(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_BO6),
.I4(CLBLM_R_X15Y141_SLICE_X21Y141_DO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y139_SLICE_X21Y139_AO5),
.O6(CLBLM_R_X15Y139_SLICE_X21Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y140_SLICE_X20Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_R_X15Y140_SLICE_X20Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y140_SLICE_X20Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_R_X15Y140_SLICE_X20Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y140_SLICE_X20Y140_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_R_X15Y140_SLICE_X20Y140_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y140_SLICE_X20Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y140_SLICE_X20Y140_DO5),
.O6(CLBLM_R_X15Y140_SLICE_X20Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y140_SLICE_X20Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y140_SLICE_X20Y140_CO5),
.O6(CLBLM_R_X15Y140_SLICE_X20Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y140_SLICE_X20Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y140_SLICE_X20Y140_BO5),
.O6(CLBLM_R_X15Y140_SLICE_X20Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y140_SLICE_X20Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y140_SLICE_X20Y140_AO5),
.O6(CLBLM_R_X15Y140_SLICE_X20Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y140_SLICE_X21Y140_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_R_X15Y140_SLICE_X21Y140_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y140_SLICE_X21Y140_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_R_X15Y140_SLICE_X21Y140_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y140_SLICE_X21Y140_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_R_X15Y140_SLICE_X21Y140_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y140_SLICE_X21Y140_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_R_X15Y140_SLICE_X21Y140_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h111111dddd11dddd)
  ) CLBLM_R_X15Y140_SLICE_X21Y140_DLUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_CO6),
.I1(CLBLM_R_X13Y139_SLICE_X19Y139_BO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I4(CLBLM_R_X15Y141_SLICE_X21Y141_BO6),
.I5(CLBLM_R_X15Y140_SLICE_X21Y140_BO6),
.O5(CLBLM_R_X15Y140_SLICE_X21Y140_DO5),
.O6(CLBLM_R_X15Y140_SLICE_X21Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0530f530053ff53f)
  ) CLBLM_R_X15Y140_SLICE_X21Y140_CLUT (
.I0(CLBLM_L_X16Y140_SLICE_X22Y140_BQ),
.I1(CLBLM_R_X15Y140_SLICE_X21Y140_CQ),
.I2(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X15Y139_SLICE_X21Y139_BQ),
.I5(CLBLM_R_X15Y140_SLICE_X20Y140_BQ),
.O5(CLBLM_R_X15Y140_SLICE_X21Y140_CO5),
.O6(CLBLM_R_X15Y140_SLICE_X21Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h227722770a0a5f5f)
  ) CLBLM_R_X15Y140_SLICE_X21Y140_BLUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I1(CLBLM_R_X15Y139_SLICE_X21Y139_AQ),
.I2(CLBLM_R_X15Y140_SLICE_X21Y140_AQ),
.I3(CLBLM_L_X16Y140_SLICE_X22Y140_AQ),
.I4(CLBLM_R_X15Y140_SLICE_X20Y140_AQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_R_X15Y140_SLICE_X21Y140_BO5),
.O6(CLBLM_R_X15Y140_SLICE_X21Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h555555550535c5f5)
  ) CLBLM_R_X15Y140_SLICE_X21Y140_ALUT (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.I1(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I2(CLBLM_R_X13Y139_SLICE_X19Y139_BO6),
.I3(CLBLM_R_X15Y141_SLICE_X21Y141_CO6),
.I4(CLBLM_R_X15Y140_SLICE_X21Y140_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y140_SLICE_X21Y140_AO5),
.O6(CLBLM_R_X15Y140_SLICE_X21Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y141_SLICE_X20Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.Q(CLBLM_R_X15Y141_SLICE_X20Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y141_SLICE_X20Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_R_X15Y141_SLICE_X20Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y141_SLICE_X20Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_R_X15Y141_SLICE_X20Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y141_SLICE_X20Y141_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_R_X15Y141_SLICE_X20Y141_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4703470347cf47cf)
  ) CLBLM_R_X15Y141_SLICE_X20Y141_DLUT (
.I0(CLBLM_R_X15Y143_SLICE_X21Y143_DO6),
.I1(CLBLM_R_X13Y139_SLICE_X19Y139_BO6),
.I2(CLBLM_R_X13Y145_SLICE_X19Y145_CO6),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I4(1'b1),
.I5(CLBLM_L_X16Y141_SLICE_X22Y141_CO6),
.O5(CLBLM_R_X15Y141_SLICE_X20Y141_DO5),
.O6(CLBLM_R_X15Y141_SLICE_X20Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLM_R_X15Y141_SLICE_X20Y141_CLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.O5(CLBLM_R_X15Y141_SLICE_X20Y141_CO5),
.O6(CLBLM_R_X15Y141_SLICE_X20Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000004000)
  ) CLBLM_R_X15Y141_SLICE_X20Y141_BLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X15Y141_SLICE_X20Y141_BO5),
.O6(CLBLM_R_X15Y141_SLICE_X20Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_R_X15Y141_SLICE_X20Y141_ALUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.O5(CLBLM_R_X15Y141_SLICE_X20Y141_AO5),
.O6(CLBLM_R_X15Y141_SLICE_X20Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y141_SLICE_X21Y141_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y139_SLICE_X21Y139_AO6),
.Q(CLBLM_R_X15Y141_SLICE_X21Y141_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y141_SLICE_X21Y141_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y141_SLICE_X21Y141_AO6),
.Q(CLBLM_R_X15Y141_SLICE_X21Y141_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y141_SLICE_X21Y141_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.Q(CLBLM_R_X15Y141_SLICE_X21Y141_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y141_SLICE_X21Y141_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_R_X15Y141_SLICE_X21Y141_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y141_SLICE_X21Y141_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y140_SLICE_X21Y140_AO6),
.Q(CLBLM_R_X15Y141_SLICE_X21Y141_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505f5f03f303f3)
  ) CLBLM_R_X15Y141_SLICE_X21Y141_DLUT (
.I0(CLBLM_L_X16Y141_SLICE_X23Y141_DQ),
.I1(CLBLM_R_X13Y141_SLICE_X19Y141_CQ),
.I2(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I3(CLBLM_R_X15Y141_SLICE_X21Y141_A5Q),
.I4(CLBLM_L_X16Y141_SLICE_X22Y141_CQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_R_X15Y141_SLICE_X21Y141_DO5),
.O6(CLBLM_R_X15Y141_SLICE_X21Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055ff550f330f33)
  ) CLBLM_R_X15Y141_SLICE_X21Y141_CLUT (
.I0(CLBLM_L_X16Y141_SLICE_X22Y141_BQ),
.I1(CLBLM_R_X15Y141_SLICE_X20Y141_DQ),
.I2(CLBLM_R_X15Y141_SLICE_X21Y141_DQ),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I4(CLBLM_L_X16Y141_SLICE_X23Y141_CQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_R_X15Y141_SLICE_X21Y141_CO5),
.O6(CLBLM_R_X15Y141_SLICE_X21Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h02138a9b4657cedf)
  ) CLBLM_R_X15Y141_SLICE_X21Y141_BLUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLM_R_X15Y141_SLICE_X21Y141_AQ),
.I3(CLBLM_R_X15Y141_SLICE_X20Y141_BQ),
.I4(CLBLM_L_X16Y141_SLICE_X23Y141_AQ),
.I5(CLBLM_R_X15Y142_SLICE_X21Y142_CQ),
.O5(CLBLM_R_X15Y141_SLICE_X21Y141_BO5),
.O6(CLBLM_R_X15Y141_SLICE_X21Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y141_SLICE_X21Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.O5(CLBLM_R_X15Y141_SLICE_X21Y141_AO5),
.O6(CLBLM_R_X15Y141_SLICE_X21Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_R_X15Y142_SLICE_X20Y142_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.Q(CLBLM_R_X15Y142_SLICE_X20Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.Q(CLBLM_R_X15Y142_SLICE_X20Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_CO6),
.Q(CLBLM_R_X15Y142_SLICE_X20Y142_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_R_X15Y142_SLICE_X20Y142_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h030303cf470347cf)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_DLUT (
.I0(CLBLM_L_X16Y142_SLICE_X22Y142_BO6),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_BO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I5(CLBLM_R_X15Y143_SLICE_X20Y143_BO6),
.O5(CLBLM_R_X15Y142_SLICE_X20Y142_DO5),
.O6(CLBLM_R_X15Y142_SLICE_X20Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.O5(CLBLM_R_X15Y142_SLICE_X20Y142_CO5),
.O6(CLBLM_R_X15Y142_SLICE_X20Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h53ff53000f0f0f0f)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_BLUT (
.I0(CLBLM_R_X15Y143_SLICE_X20Y143_CO6),
.I1(CLBLM_L_X16Y142_SLICE_X22Y142_DO6),
.I2(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_BO6),
.I4(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y142_SLICE_X20Y142_BO5),
.O6(CLBLM_R_X15Y142_SLICE_X20Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555533550f55)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_ALUT (
.I0(CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O),
.I1(CLBLM_R_X15Y142_SLICE_X21Y142_DO6),
.I2(CLBLM_R_X15Y142_SLICE_X21Y142_CO6),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_BO6),
.I4(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I5(1'b1),
.O5(CLBLM_R_X15Y142_SLICE_X20Y142_AO5),
.O6(CLBLM_R_X15Y142_SLICE_X20Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_R_X15Y142_SLICE_X21Y142_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X21Y142_AO6),
.Q(CLBLM_R_X15Y142_SLICE_X21Y142_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.Q(CLBLM_R_X15Y142_SLICE_X21Y142_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_L_X16Y136_SLICE_X22Y136_AO6),
.Q(CLBLM_R_X15Y142_SLICE_X21Y142_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y141_SLICE_X22Y141_BO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.Q(CLBLM_R_X15Y142_SLICE_X21Y142_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033ccff47474747)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_DLUT (
.I0(CLBLM_R_X15Y140_SLICE_X21Y140_BQ),
.I1(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I2(CLBLM_R_X15Y143_SLICE_X21Y143_B5Q),
.I3(CLBLM_L_X16Y143_SLICE_X22Y143_CQ),
.I4(CLBLM_R_X15Y142_SLICE_X20Y142_C5Q),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_R_X15Y142_SLICE_X21Y142_DO5),
.O6(CLBLM_R_X15Y142_SLICE_X21Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00331d1dccff1d1d)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_CLUT (
.I0(CLBLM_R_X13Y141_SLICE_X19Y141_BQ),
.I1(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I2(CLBLM_R_X15Y144_SLICE_X21Y144_CQ),
.I3(CLBLM_R_X15Y142_SLICE_X21Y142_A5Q),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(CLBLM_L_X16Y142_SLICE_X22Y142_DQ),
.O5(CLBLM_R_X15Y142_SLICE_X21Y142_CO5),
.O6(CLBLM_R_X15Y142_SLICE_X21Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h111105afbbbb05af)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_BLUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I1(CLBLM_R_X15Y142_SLICE_X21Y142_BQ),
.I2(CLBLM_R_X15Y141_SLICE_X20Y141_AQ),
.I3(CLBLM_R_X15Y144_SLICE_X21Y144_BQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I5(CLBLM_L_X16Y142_SLICE_X22Y142_BQ),
.O5(CLBLM_R_X15Y142_SLICE_X21Y142_BO5),
.O6(CLBLM_R_X15Y142_SLICE_X21Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.O5(CLBLM_R_X15Y142_SLICE_X21Y142_AO5),
.O6(CLBLM_R_X15Y142_SLICE_X21Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y143_SLICE_X20Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.Q(CLBLM_R_X15Y143_SLICE_X20Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y143_SLICE_X20Y143_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.Q(CLBLM_R_X15Y143_SLICE_X20Y143_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y143_SLICE_X20Y143_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.Q(CLBLM_R_X15Y143_SLICE_X20Y143_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y143_SLICE_X20Y143_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_R_X15Y143_SLICE_X20Y143_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a5f5f22772277)
  ) CLBLM_R_X15Y143_SLICE_X20Y143_DLUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I1(CLBLM_R_X15Y143_SLICE_X20Y143_CQ),
.I2(CLBLM_R_X15Y142_SLICE_X20Y142_CQ),
.I3(CLBLM_R_X15Y143_SLICE_X21Y143_CQ),
.I4(CLBLM_R_X15Y144_SLICE_X20Y144_CQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_R_X15Y143_SLICE_X20Y143_DO5),
.O6(CLBLM_R_X15Y143_SLICE_X20Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0035f0350f35ff35)
  ) CLBLM_R_X15Y143_SLICE_X20Y143_CLUT (
.I0(CLBLM_R_X15Y143_SLICE_X21Y143_AQ),
.I1(CLBLM_R_X15Y143_SLICE_X20Y143_AQ),
.I2(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X15Y142_SLICE_X20Y142_AQ),
.I5(CLBLM_R_X15Y144_SLICE_X20Y144_BQ),
.O5(CLBLM_R_X15Y143_SLICE_X20Y143_CO5),
.O6(CLBLM_R_X15Y143_SLICE_X20Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800bb00c000f300)
  ) CLBLM_R_X15Y143_SLICE_X20Y143_BLUT (
.I0(CLBLM_R_X15Y142_SLICE_X20Y142_AQ),
.I1(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I2(CLBLM_R_X15Y143_SLICE_X20Y143_AQ),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I4(CLBLM_R_X15Y143_SLICE_X20Y143_AO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_R_X15Y143_SLICE_X20Y143_BO5),
.O6(CLBLM_R_X15Y143_SLICE_X20Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h330033ff00550055)
  ) CLBLM_R_X15Y143_SLICE_X20Y143_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.I1(CLBLM_R_X15Y144_SLICE_X20Y144_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I4(CLBLM_R_X15Y143_SLICE_X21Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y143_SLICE_X20Y143_AO5),
.O6(CLBLM_R_X15Y143_SLICE_X20Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y143_SLICE_X21Y143_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_R_X15Y143_SLICE_X21Y143_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y143_SLICE_X21Y143_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.Q(CLBLM_R_X15Y143_SLICE_X21Y143_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y143_SLICE_X21Y143_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_BO6),
.Q(CLBLM_R_X15Y143_SLICE_X21Y143_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y143_SLICE_X21Y143_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.Q(CLBLM_R_X15Y143_SLICE_X21Y143_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y143_SLICE_X21Y143_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_R_X15Y143_SLICE_X21Y143_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33553355000fff0f)
  ) CLBLM_R_X15Y143_SLICE_X21Y143_DLUT (
.I0(CLBLM_L_X16Y143_SLICE_X22Y143_BQ),
.I1(CLBLM_R_X15Y142_SLICE_X20Y142_DQ),
.I2(CLBLM_R_X15Y143_SLICE_X21Y143_DQ),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I4(CLBLM_R_X15Y143_SLICE_X20Y143_DQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.O5(CLBLM_R_X15Y143_SLICE_X21Y143_DO5),
.O6(CLBLM_R_X15Y143_SLICE_X21Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc474733ff4747)
  ) CLBLM_R_X15Y143_SLICE_X21Y143_CLUT (
.I0(CLBLM_L_X16Y143_SLICE_X22Y143_AQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.I2(CLBLM_R_X15Y143_SLICE_X21Y143_BQ),
.I3(CLBLM_R_X15Y142_SLICE_X20Y142_BQ),
.I4(CLBLM_R_X13Y139_SLICE_X19Y139_DO6),
.I5(CLBLM_R_X15Y143_SLICE_X20Y143_BQ),
.O5(CLBLM_R_X15Y143_SLICE_X21Y143_CO5),
.O6(CLBLM_R_X15Y143_SLICE_X21Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000000)
  ) CLBLM_R_X15Y143_SLICE_X21Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.O5(CLBLM_R_X15Y143_SLICE_X21Y143_BO5),
.O6(CLBLM_R_X15Y143_SLICE_X21Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0533af3333333333)
  ) CLBLM_R_X15Y143_SLICE_X21Y143_ALUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.I1(CLBLM_R_X15Y144_SLICE_X21Y144_AO6),
.I2(CLBLM_R_X15Y142_SLICE_X21Y142_BO6),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_BO6),
.I4(CLBLM_R_X15Y143_SLICE_X21Y143_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.O6(CLBLM_R_X15Y143_SLICE_X21Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y143_SLICE_X22Y143_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.Q(CLBLM_R_X15Y144_SLICE_X20Y144_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_L_X16Y143_SLICE_X22Y143_AO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y144_SLICE_X21Y144_BO6),
.Q(CLBLM_R_X15Y144_SLICE_X20Y144_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y144_SLICE_X20Y144_DO5),
.O6(CLBLM_R_X15Y144_SLICE_X20Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haffa0faa30af3f50)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_CLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_AO6),
.I2(CLBLM_R_X15Y146_SLICE_X20Y146_AO6),
.I3(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.O5(CLBLM_R_X15Y144_SLICE_X20Y144_CO5),
.O6(CLBLM_R_X15Y144_SLICE_X20Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffffbb0088)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I5(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.O5(CLBLM_R_X15Y144_SLICE_X20Y144_BO5),
.O6(CLBLM_R_X15Y144_SLICE_X20Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a0fffaa5faa5)
  ) CLBLM_R_X15Y144_SLICE_X20Y144_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I4(CLBLM_R_X13Y144_SLICE_X19Y144_CO5),
.I5(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.O5(CLBLM_R_X15Y144_SLICE_X20Y144_AO5),
.O6(CLBLM_R_X15Y144_SLICE_X20Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X15Y144_SLICE_X20Y144_MUXF7A (
.I0(CLBLM_R_X15Y144_SLICE_X20Y144_BO6),
.I1(CLBLM_R_X15Y144_SLICE_X20Y144_AO6),
.O(CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O),
.S(CLBLM_R_X15Y146_SLICE_X20Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y145_SLICE_X20Y145_CO6),
.Q(CLBLM_R_X15Y144_SLICE_X21Y144_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y143_SLICE_X21Y143_AO5),
.Q(CLBLM_R_X15Y144_SLICE_X21Y144_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(CLBLM_R_X15Y141_SLICE_X20Y141_CO6),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_R_X15Y144_SLICE_X21Y144_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y144_SLICE_X21Y144_DO5),
.O6(CLBLM_R_X15Y144_SLICE_X21Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcffc0fcc50cf5f30)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_CLUT (
.I0(CLBLM_L_X12Y144_SLICE_X17Y144_CO6),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I2(CLBLM_R_X15Y146_SLICE_X20Y146_AO6),
.I3(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.O5(CLBLM_R_X15Y144_SLICE_X21Y144_CO5),
.O6(CLBLM_R_X15Y144_SLICE_X21Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2afa2a50132d132d)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_BLUT (
.I0(CLBLM_R_X15Y146_SLICE_X20Y146_AO6),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I4(CLBLM_L_X12Y144_SLICE_X17Y144_CO6),
.I5(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.O5(CLBLM_R_X15Y144_SLICE_X21Y144_BO5),
.O6(CLBLM_R_X15Y144_SLICE_X21Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88f0ff33ee99aacc)
  ) CLBLM_R_X15Y144_SLICE_X21Y144_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I2(CLBLM_R_X13Y144_SLICE_X19Y144_CO6),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I4(CLBLM_R_X15Y146_SLICE_X20Y146_AO6),
.I5(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.O5(CLBLM_R_X15Y144_SLICE_X21Y144_AO5),
.O6(CLBLM_R_X15Y144_SLICE_X21Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y145_SLICE_X20Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y145_SLICE_X20Y145_DO5),
.O6(CLBLM_R_X15Y145_SLICE_X20Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a00af55a5a5f0a5)
  ) CLBLM_R_X15Y145_SLICE_X20Y145_CLUT (
.I0(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I3(CLBLM_R_X15Y146_SLICE_X20Y146_AO6),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.O5(CLBLM_R_X15Y145_SLICE_X20Y145_CO5),
.O6(CLBLM_R_X15Y145_SLICE_X20Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcff0cff0cfb8cfb8)
  ) CLBLM_R_X15Y145_SLICE_X20Y145_BLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I3(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.O5(CLBLM_R_X15Y145_SLICE_X20Y145_BO5),
.O6(CLBLM_R_X15Y145_SLICE_X20Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80b380b3e9e9e9e9)
  ) CLBLM_R_X15Y145_SLICE_X20Y145_ALUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I3(CLBLM_R_X13Y145_SLICE_X19Y145_BO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y146_SLICE_X19Y146_AO6),
.O5(CLBLM_R_X15Y145_SLICE_X20Y145_AO5),
.O6(CLBLM_R_X15Y145_SLICE_X20Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X15Y145_SLICE_X20Y145_MUXF7A (
.I0(CLBLM_R_X15Y145_SLICE_X20Y145_BO6),
.I1(CLBLM_R_X15Y145_SLICE_X20Y145_AO6),
.O(CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O),
.S(CLBLM_R_X15Y146_SLICE_X20Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y145_SLICE_X21Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y145_SLICE_X21Y145_DO5),
.O6(CLBLM_R_X15Y145_SLICE_X21Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y145_SLICE_X21Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y145_SLICE_X21Y145_CO5),
.O6(CLBLM_R_X15Y145_SLICE_X21Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y145_SLICE_X21Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y145_SLICE_X21Y145_BO5),
.O6(CLBLM_R_X15Y145_SLICE_X21Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y145_SLICE_X21Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y145_SLICE_X21Y145_AO5),
.O6(CLBLM_R_X15Y145_SLICE_X21Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y146_SLICE_X20Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y146_SLICE_X20Y146_DO5),
.O6(CLBLM_R_X15Y146_SLICE_X20Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y146_SLICE_X20Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y146_SLICE_X20Y146_CO5),
.O6(CLBLM_R_X15Y146_SLICE_X20Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y146_SLICE_X20Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y146_SLICE_X20Y146_BO5),
.O6(CLBLM_R_X15Y146_SLICE_X20Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050a000a0500000)
  ) CLBLM_R_X15Y146_SLICE_X20Y146_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.O5(CLBLM_R_X15Y146_SLICE_X20Y146_AO5),
.O6(CLBLM_R_X15Y146_SLICE_X20Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h02a057ff0200575f)
  ) CLBLM_R_X15Y146_SLICE_X21Y146_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I5(CLBLM_R_X13Y145_SLICE_X19Y145_BO6),
.O5(CLBLM_R_X15Y146_SLICE_X21Y146_DO5),
.O6(CLBLM_R_X15Y146_SLICE_X21Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8fa50f0f0f0f0)
  ) CLBLM_R_X15Y146_SLICE_X21Y146_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I3(CLBLM_R_X13Y144_SLICE_X19Y144_CO6),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.O5(CLBLM_R_X15Y146_SLICE_X21Y146_CO5),
.O6(CLBLM_R_X15Y146_SLICE_X21Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0555f5550aeafaea)
  ) CLBLM_R_X15Y146_SLICE_X21Y146_BLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.O5(CLBLM_R_X15Y146_SLICE_X21Y146_BO5),
.O6(CLBLM_R_X15Y146_SLICE_X21Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeeaaaeaaaeaa)
  ) CLBLM_R_X15Y146_SLICE_X21Y146_ALUT (
.I0(CLBLM_R_X15Y146_SLICE_X21Y146_DO6),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.O5(CLBLM_R_X15Y146_SLICE_X21Y146_AO5),
.O6(CLBLM_R_X15Y146_SLICE_X21Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_R_X15Y146_SLICE_X21Y146_MUXF7A (
.I0(CLBLM_R_X15Y146_SLICE_X21Y146_BO6),
.I1(CLBLM_R_X15Y146_SLICE_X21Y146_AO6),
.O(CLBLM_R_X15Y146_SLICE_X21Y146_F7AMUX_O),
.S(CLBLM_R_X15Y150_SLICE_X20Y150_DO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y147_SLICE_X20Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y147_SLICE_X20Y147_DO5),
.O6(CLBLM_R_X15Y147_SLICE_X20Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y147_SLICE_X20Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y147_SLICE_X20Y147_CO5),
.O6(CLBLM_R_X15Y147_SLICE_X20Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y147_SLICE_X20Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y147_SLICE_X20Y147_BO5),
.O6(CLBLM_R_X15Y147_SLICE_X20Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y147_SLICE_X20Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y147_SLICE_X20Y147_AO5),
.O6(CLBLM_R_X15Y147_SLICE_X20Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y147_SLICE_X21Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y147_SLICE_X21Y147_DO5),
.O6(CLBLM_R_X15Y147_SLICE_X21Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y147_SLICE_X21Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y147_SLICE_X21Y147_CO5),
.O6(CLBLM_R_X15Y147_SLICE_X21Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y147_SLICE_X21Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y147_SLICE_X21Y147_BO5),
.O6(CLBLM_R_X15Y147_SLICE_X21Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50005fff5fff50c0)
  ) CLBLM_R_X15Y147_SLICE_X21Y147_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.O5(CLBLM_R_X15Y147_SLICE_X21Y147_AO5),
.O6(CLBLM_R_X15Y147_SLICE_X21Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y148_SLICE_X20Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y148_SLICE_X20Y148_DO5),
.O6(CLBLM_R_X15Y148_SLICE_X20Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff88a2ffffffff)
  ) CLBLM_R_X15Y148_SLICE_X20Y148_CLUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I5(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.O5(CLBLM_R_X15Y148_SLICE_X20Y148_CO5),
.O6(CLBLM_R_X15Y148_SLICE_X20Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7000ffff8080)
  ) CLBLM_R_X15Y148_SLICE_X20Y148_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I3(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.O5(CLBLM_R_X15Y148_SLICE_X20Y148_BO5),
.O6(CLBLM_R_X15Y148_SLICE_X20Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaafeae)
  ) CLBLM_R_X15Y148_SLICE_X20Y148_ALUT (
.I0(CLBLM_R_X15Y148_SLICE_X20Y148_BO6),
.I1(CLBLM_R_X15Y150_SLICE_X21Y150_CO6),
.I2(CLBLM_R_X15Y152_SLICE_X20Y152_DO6),
.I3(CLBLM_L_X16Y152_SLICE_X22Y152_D_XOR),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(CLBLM_R_X15Y148_SLICE_X20Y148_CO6),
.O5(CLBLM_R_X15Y148_SLICE_X20Y148_AO5),
.O6(CLBLM_R_X15Y148_SLICE_X20Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h56006a00a9ff95ff)
  ) CLBLM_R_X15Y148_SLICE_X21Y148_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.O5(CLBLM_R_X15Y148_SLICE_X21Y148_DO5),
.O6(CLBLM_R_X15Y148_SLICE_X21Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdf80805fff00a0)
  ) CLBLM_R_X15Y148_SLICE_X21Y148_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_R_X15Y148_SLICE_X21Y148_AO5),
.I4(CLBLM_R_X15Y148_SLICE_X21Y148_DO6),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.O5(CLBLM_R_X15Y148_SLICE_X21Y148_CO5),
.O6(CLBLM_R_X15Y148_SLICE_X21Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0faaccff0faacc00)
  ) CLBLM_R_X15Y148_SLICE_X21Y148_BLUT (
.I0(CLBLM_R_X15Y147_SLICE_X21Y147_AO6),
.I1(CLBLM_R_X15Y149_SLICE_X21Y149_AO6),
.I2(CLBLM_R_X15Y146_SLICE_X21Y146_CO6),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I5(CLBLM_R_X15Y148_SLICE_X21Y148_CO6),
.O5(CLBLM_R_X15Y148_SLICE_X21Y148_BO5),
.O6(CLBLM_R_X15Y148_SLICE_X21Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69696969b24d4db2)
  ) CLBLM_R_X15Y148_SLICE_X21Y148_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y148_SLICE_X21Y148_AO5),
.O6(CLBLM_R_X15Y148_SLICE_X21Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff00ff)
  ) CLBLM_R_X15Y149_SLICE_X20Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.O5(CLBLM_R_X15Y149_SLICE_X20Y149_DO5),
.O6(CLBLM_R_X15Y149_SLICE_X20Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff55f555d7)
  ) CLBLM_R_X15Y149_SLICE_X20Y149_CLUT (
.I0(CLBLM_R_X15Y149_SLICE_X20Y149_AO6),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.I4(CLBLM_R_X15Y149_SLICE_X20Y149_BO5),
.I5(CLBLM_R_X13Y149_SLICE_X19Y149_AO6),
.O5(CLBLM_R_X15Y149_SLICE_X20Y149_CO5),
.O6(CLBLM_R_X15Y149_SLICE_X20Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c400c4c4c40000)
  ) CLBLM_R_X15Y149_SLICE_X20Y149_BLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(CLBLM_R_X13Y149_SLICE_X19Y149_AO6),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y149_SLICE_X20Y149_BO5),
.O6(CLBLM_R_X15Y149_SLICE_X20Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0000bfbfffff)
  ) CLBLM_R_X15Y149_SLICE_X20Y149_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y149_SLICE_X20Y149_AO5),
.O6(CLBLM_R_X15Y149_SLICE_X20Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y149_SLICE_X21Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y149_SLICE_X21Y149_DO5),
.O6(CLBLM_R_X15Y149_SLICE_X21Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y149_SLICE_X21Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y149_SLICE_X21Y149_CO5),
.O6(CLBLM_R_X15Y149_SLICE_X21Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y149_SLICE_X21Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y149_SLICE_X21Y149_BO5),
.O6(CLBLM_R_X15Y149_SLICE_X21Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f500f500cfcfc0c)
  ) CLBLM_R_X15Y149_SLICE_X21Y149_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I1(CLBLM_R_X15Y152_SLICE_X21Y152_BO6),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.I4(CLBLM_R_X15Y149_SLICE_X20Y149_DO6),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.O5(CLBLM_R_X15Y149_SLICE_X21Y149_AO5),
.O6(CLBLM_R_X15Y149_SLICE_X21Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y150_SLICE_X20Y150_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y150_SLICE_X20Y150_AO6),
.Q(CLBLM_R_X15Y150_SLICE_X20Y150_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLM_R_X15Y150_SLICE_X20Y150_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.O6(CLBLM_R_X15Y150_SLICE_X20Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2800220082008800)
  ) CLBLM_R_X15Y150_SLICE_X20Y150_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.I5(CLBLM_R_X13Y149_SLICE_X19Y149_AO6),
.O5(CLBLM_R_X15Y150_SLICE_X20Y150_CO5),
.O6(CLBLM_R_X15Y150_SLICE_X20Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcbcb0000cbcbccff)
  ) CLBLM_R_X15Y150_SLICE_X20Y150_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I3(CLBLM_R_X15Y152_SLICE_X20Y152_BO6),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I5(CLBLM_R_X15Y150_SLICE_X20Y150_CO6),
.O5(CLBLM_R_X15Y150_SLICE_X20Y150_BO5),
.O6(CLBLM_R_X15Y150_SLICE_X20Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e1f0f0f0f0f0f0)
  ) CLBLM_R_X15Y150_SLICE_X20Y150_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.O5(CLBLM_R_X15Y150_SLICE_X20Y150_AO5),
.O6(CLBLM_R_X15Y150_SLICE_X20Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0d0d0d0a0f5a0f5)
  ) CLBLM_R_X15Y150_SLICE_X21Y150_DLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_A5Q),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(1'b1),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_R_X15Y150_SLICE_X21Y150_DO5),
.O6(CLBLM_R_X15Y150_SLICE_X21Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefff0100ef0001)
  ) CLBLM_R_X15Y150_SLICE_X21Y150_CLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I3(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I4(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.I5(CLBLM_L_X16Y150_SLICE_X22Y150_C_XOR),
.O5(CLBLM_R_X15Y150_SLICE_X21Y150_CO5),
.O6(CLBLM_R_X15Y150_SLICE_X21Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1aaf1aa015af15a0)
  ) CLBLM_R_X15Y150_SLICE_X21Y150_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I4(CLBLM_L_X16Y152_SLICE_X23Y152_BO6),
.I5(CLBLM_R_X15Y149_SLICE_X20Y149_BO6),
.O5(CLBLM_R_X15Y150_SLICE_X21Y150_BO5),
.O6(CLBLM_R_X15Y150_SLICE_X21Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0ff00dd11)
  ) CLBLM_R_X15Y150_SLICE_X21Y150_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I1(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_A5Q),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y150_SLICE_X21Y150_AO5),
.O6(CLBLM_R_X15Y150_SLICE_X21Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y151_SLICE_X20Y151_CO6),
.Q(CLBLM_R_X15Y151_SLICE_X20Y151_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y151_SLICE_X20Y151_CO5),
.Q(CLBLM_R_X15Y151_SLICE_X20Y151_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he0e0eee0a0a0aaa0)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_DLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I3(CLBLM_R_X15Y151_SLICE_X20Y151_AO5),
.I4(CLBLM_R_X15Y151_SLICE_X20Y151_BO5),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_DO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccff00f0f0)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_CLUT (
.I0(CLBLM_L_X16Y152_SLICE_X22Y152_D_XOR),
.I1(CLBLM_R_X15Y150_SLICE_X21Y150_CO6),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_BO6),
.I3(CLBLM_L_X16Y153_SLICE_X22Y153_D_XOR),
.I4(CLBLM_R_X15Y152_SLICE_X20Y152_DO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_CO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003333757f757f)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_BO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffaf00a000)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_AO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_A5_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y152_SLICE_X21Y152_CO6),
.Q(CLBLM_R_X15Y151_SLICE_X21Y151_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y151_SLICE_X21Y151_AO6),
.Q(CLBLM_R_X15Y151_SLICE_X21Y151_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafcfa0cfafc0a0c0)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_DO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddf588f5dda088a0)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_CLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_CO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fdcd3101)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_BLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I1(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I2(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I3(CLBLM_R_X15Y151_SLICE_X20Y151_BQ),
.I4(CLBLM_L_X16Y151_SLICE_X22Y151_C_XOR),
.I5(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_BO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0e1f0f0f0)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I1(CLBLM_R_X15Y150_SLICE_X20Y150_DO6),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I3(CLBLM_R_X15Y150_SLICE_X20Y150_DO5),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_AO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y152_SLICE_X20Y152_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y152_SLICE_X20Y152_BO6),
.Q(CLBLM_R_X15Y152_SLICE_X20Y152_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_R_X15Y152_SLICE_X20Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X15Y151_SLICE_X20Y151_DO6),
.I4(1'b1),
.I5(CLBLM_L_X16Y154_SLICE_X22Y154_A_CY),
.O5(CLBLM_R_X15Y152_SLICE_X20Y152_DO5),
.O6(CLBLM_R_X15Y152_SLICE_X20Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c8c8c8cdcdcdcd)
  ) CLBLM_R_X15Y152_SLICE_X20Y152_CLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(CLBLM_R_X15Y152_SLICE_X20Y152_AQ),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.O5(CLBLM_R_X15Y152_SLICE_X20Y152_CO5),
.O6(CLBLM_R_X15Y152_SLICE_X20Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bbbbbb888888)
  ) CLBLM_R_X15Y152_SLICE_X20Y152_BLUT (
.I0(CLBLM_L_X16Y153_SLICE_X22Y153_B_XOR),
.I1(CLBLM_R_X15Y152_SLICE_X20Y152_DO6),
.I2(1'b1),
.I3(CLBLM_L_X16Y151_SLICE_X22Y151_A_XOR),
.I4(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I5(CLBLM_R_X15Y152_SLICE_X20Y152_CO6),
.O5(CLBLM_R_X15Y152_SLICE_X20Y152_BO5),
.O6(CLBLM_R_X15Y152_SLICE_X20Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcecfd30302031)
  ) CLBLM_R_X15Y152_SLICE_X20Y152_ALUT (
.I0(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I1(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I2(CLBLM_R_X15Y152_SLICE_X20Y152_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I5(CLBLM_L_X16Y151_SLICE_X22Y151_A_XOR),
.O5(CLBLM_R_X15Y152_SLICE_X20Y152_AO5),
.O6(CLBLM_R_X15Y152_SLICE_X20Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y152_SLICE_X21Y152_A_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y152_SLICE_X21Y152_BO6),
.Q(CLBLM_R_X15Y152_SLICE_X21Y152_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y152_SLICE_X21Y152_B_FDCE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.CLR(LIOB33_X0Y105_IOB_X0Y106_I),
.D(CLBLM_R_X15Y153_SLICE_X21Y153_CO6),
.Q(CLBLM_R_X15Y152_SLICE_X21Y152_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa0000ffff0055)
  ) CLBLM_R_X15Y152_SLICE_X21Y152_DLUT (
.I0(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I4(CLBLM_R_X15Y152_SLICE_X21Y152_AQ),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.O5(CLBLM_R_X15Y152_SLICE_X21Y152_DO5),
.O6(CLBLM_R_X15Y152_SLICE_X21Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefef4f40e0e0404)
  ) CLBLM_R_X15Y152_SLICE_X21Y152_CLUT (
.I0(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I1(CLBLM_R_X15Y150_SLICE_X21Y150_AO5),
.I2(CLBLM_R_X15Y152_SLICE_X20Y152_DO6),
.I3(1'b1),
.I4(CLBLM_L_X16Y150_SLICE_X22Y150_B_XOR),
.I5(CLBLM_L_X16Y152_SLICE_X22Y152_C_XOR),
.O5(CLBLM_R_X15Y152_SLICE_X21Y152_CO5),
.O6(CLBLM_R_X15Y152_SLICE_X21Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffccaaaa3300)
  ) CLBLM_R_X15Y152_SLICE_X21Y152_BLUT (
.I0(CLBLM_L_X16Y152_SLICE_X22Y152_B_XOR),
.I1(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I2(1'b1),
.I3(CLBLM_R_X15Y152_SLICE_X21Y152_DO6),
.I4(CLBLM_R_X15Y152_SLICE_X20Y152_DO6),
.I5(CLBLM_L_X16Y150_SLICE_X22Y150_A_XOR),
.O5(CLBLM_R_X15Y152_SLICE_X21Y152_BO5),
.O6(CLBLM_R_X15Y152_SLICE_X21Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbbff00008800)
  ) CLBLM_R_X15Y152_SLICE_X21Y152_ALUT (
.I0(CLBLM_L_X16Y150_SLICE_X22Y150_B_XOR),
.I1(CLBLM_R_X15Y151_SLICE_X20Y151_DO6),
.I2(1'b1),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_DO6),
.I4(CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR),
.I5(CLBLM_R_X15Y150_SLICE_X21Y150_AO5),
.O5(CLBLM_R_X15Y152_SLICE_X21Y152_AO5),
.O6(CLBLM_R_X15Y152_SLICE_X21Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X20Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X20Y153_DO5),
.O6(CLBLM_R_X15Y153_SLICE_X20Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X20Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X20Y153_CO5),
.O6(CLBLM_R_X15Y153_SLICE_X20Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X20Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X20Y153_BO5),
.O6(CLBLM_R_X15Y153_SLICE_X20Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X20Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X20Y153_AO5),
.O6(CLBLM_R_X15Y153_SLICE_X20Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X21Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X21Y153_DO5),
.O6(CLBLM_R_X15Y153_SLICE_X21Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfc0c0c0cfc0)
  ) CLBLM_R_X15Y153_SLICE_X21Y153_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X16Y153_SLICE_X22Y153_A_XOR),
.I2(CLBLM_R_X15Y152_SLICE_X20Y152_DO6),
.I3(CLBLM_R_X15Y153_SLICE_X21Y153_AO5),
.I4(CLBLM_L_X16Y153_SLICE_X23Y153_AO6),
.I5(CLBLM_L_X16Y150_SLICE_X22Y150_D_XOR),
.O5(CLBLM_R_X15Y153_SLICE_X21Y153_CO5),
.O6(CLBLM_R_X15Y153_SLICE_X21Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcffffff0c000000)
  ) CLBLM_R_X15Y153_SLICE_X21Y153_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X16Y150_SLICE_X22Y150_D_XOR),
.I2(CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR),
.I3(CLBLM_R_X15Y151_SLICE_X21Y151_DO6),
.I4(CLBLM_R_X15Y151_SLICE_X20Y151_DO6),
.I5(CLBLM_R_X15Y153_SLICE_X21Y153_AO5),
.O5(CLBLM_R_X15Y153_SLICE_X21Y153_BO5),
.O6(CLBLM_R_X15Y153_SLICE_X21Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0ccccc0cf)
  ) CLBLM_R_X15Y153_SLICE_X21Y153_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X15Y152_SLICE_X21Y152_BQ),
.I2(CLBLM_R_X15Y151_SLICE_X21Y151_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I4(CLBLM_R_X15Y150_SLICE_X20Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X21Y153_AO5),
.O6(CLBLM_R_X15Y153_SLICE_X21Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y51_IOB_X0Y51_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.O(LIOB33_X0Y51_IOB_X0Y51_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y51_IOB_X0Y52_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.O(LIOB33_X0Y51_IOB_X0Y52_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y53_IOB_X0Y53_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X5Y135_B5Q),
.O(LIOB33_X0Y53_IOB_X0Y53_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y53_IOB_X0Y54_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.O(LIOB33_X0Y53_IOB_X0Y54_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y55_IOB_X0Y55_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.O(LIOB33_X0Y55_IOB_X0Y55_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y55_IOB_X0Y56_OBUF (
.I(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.O(LIOB33_X0Y55_IOB_X0Y56_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y57_IOB_X0Y57_OBUF (
.I(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.O(LIOB33_X0Y57_IOB_X0Y57_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y57_IOB_X0Y58_OBUF (
.I(CLBLM_R_X5Y136_SLICE_X7Y136_DQ),
.O(LIOB33_X0Y57_IOB_X0Y58_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y59_IOB_X0Y59_OBUF (
.I(CLBLM_L_X12Y128_SLICE_X16Y128_AQ),
.O(LIOB33_X0Y59_IOB_X0Y59_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y59_IOB_X0Y60_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.O(LIOB33_X0Y59_IOB_X0Y60_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y61_IOB_X0Y61_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.O(LIOB33_X0Y61_IOB_X0Y61_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y61_IOB_X0Y62_OBUF (
.I(CLBLL_L_X2Y116_SLICE_X0Y116_AQ),
.O(LIOB33_X0Y61_IOB_X0Y62_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y63_OBUF (
.I(1'b1),
.O(LIOB33_X0Y63_IOB_X0Y63_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X4Y135_B5Q),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X4Y135_C5Q),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X4Y135_DQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X1Y135_AQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLL_L_X2Y135_SLICE_X1Y135_A5Q),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X5Y135_A5Q),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y138_SLICE_X1Y138_AO6),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X2Y137_SLICE_X0Y137_AO6),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLL_L_X2Y137_SLICE_X0Y137_AO5),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X2Y137_SLICE_X1Y137_AO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X2Y137_SLICE_X1Y137_AO5),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X2Y137_SLICE_X1Y137_BO6),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X2Y137_SLICE_X1Y137_BO5),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X1Y139_DO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X1Y139_DO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X1Y139_AO6),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X1Y139_AO5),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X1Y139_BO6),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X1Y139_BO5),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X1Y139_CO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X1Y139_CO5),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X2Y143_SLICE_X0Y143_AQ),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X2Y144_SLICE_X0Y144_AQ),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X2Y144_SLICE_X0Y144_A5Q),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLL_L_X2Y145_SLICE_X0Y145_AQ),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_L_X2Y145_SLICE_X0Y145_A5Q),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X2Y147_SLICE_X0Y147_AQ),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y151_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y151_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y152_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y152_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y153_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y153_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y154_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y154_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y155_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y156_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y156_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y157_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y157_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y158_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y158_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y159_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y159_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y160_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y160_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y161_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y161_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y162_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y162_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y163_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y163_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y164_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y164_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y165_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y165_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y166_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y166_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y167_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y167_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y168_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y168_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y169_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y169_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y170_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y170_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y171_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y171_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y172_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y172_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y173_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y173_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y173_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y174_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y174_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y174_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y175_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y175_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y175_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y176_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y176_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y176_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y177_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y177_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y177_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y178_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y178_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y178_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y179_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y179_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y179_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y180_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y180_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y180_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y181_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y181_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y181_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y182_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y182_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y182_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y183_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y183_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y183_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y184_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y184_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y184_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y185_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y185_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y185_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y186_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y186_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y186_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y187_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y187_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y187_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y188_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y188_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y188_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y189_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y189_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y189_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y190_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y190_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y190_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y191_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y191_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y191_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y192_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y192_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y192_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y193_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y193_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y193_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y194_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y194_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y194_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y195_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y195_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y195_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y196_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y196_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y196_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y197_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y197_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y197_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y198_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y198_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y198_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y50_IOB_X0Y50_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLL_L_X2Y147_SLICE_X0Y147_A5Q),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y150_IOB_X0Y150_IBUF (
.I(LIOB33_SING_X0Y150_IOB_X0Y150_IPAD),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y199_IOB_X0Y199_IBUF (
.I(LIOB33_SING_X0Y199_IOB_X0Y199_IPAD),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y124_OBUF (
.I(CLBLM_L_X16Y133_SLICE_X23Y133_AQ),
.O(RIOB33_X105Y123_IOB_X1Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y125_OBUF (
.I(CLBLM_L_X16Y133_SLICE_X22Y133_AQ),
.O(RIOB33_X105Y125_IOB_X1Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y126_OBUF (
.I(CLBLM_L_X16Y133_SLICE_X23Y133_BQ),
.O(RIOB33_X105Y125_IOB_X1Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(CLBLM_L_X16Y133_SLICE_X22Y133_BQ),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(CLBLM_L_X16Y133_SLICE_X23Y133_CQ),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(CLBLM_L_X16Y134_SLICE_X23Y134_AQ),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(CLBLM_L_X16Y133_SLICE_X23Y133_DQ),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(CLBLM_L_X16Y133_SLICE_X22Y133_CQ),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(CLBLM_L_X16Y135_SLICE_X22Y135_AQ),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(CLBLM_L_X16Y134_SLICE_X22Y134_BQ),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(CLBLM_L_X16Y135_SLICE_X23Y135_AQ),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(CLBLM_L_X16Y135_SLICE_X22Y135_BQ),
.O(RIOB33_X105Y135_IOB_X1Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(CLBLM_L_X16Y136_SLICE_X23Y136_BQ),
.O(RIOB33_X105Y137_IOB_X1Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(CLBLM_L_X16Y136_SLICE_X23Y136_CQ),
.O(RIOB33_X105Y137_IOB_X1Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(CLBLM_L_X16Y138_SLICE_X23Y138_AQ),
.O(RIOB33_X105Y139_IOB_X1Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(CLBLM_L_X16Y139_SLICE_X22Y139_AQ),
.O(RIOB33_X105Y139_IOB_X1Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(CLBLM_R_X13Y138_SLICE_X19Y138_AQ),
.O(RIOB33_X105Y141_IOB_X1Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(CLBLM_R_X13Y138_SLICE_X19Y138_BQ),
.O(RIOB33_X105Y141_IOB_X1Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(CLBLM_L_X16Y136_SLICE_X23Y136_DQ),
.O(RIOB33_X105Y143_IOB_X1Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(CLBLM_R_X13Y138_SLICE_X19Y138_CQ),
.O(RIOB33_X105Y143_IOB_X1Y144_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(CLBLM_L_X16Y138_SLICE_X22Y138_AQ),
.O(RIOB33_X105Y145_IOB_X1Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y146_OBUF (
.I(CLBLM_L_X16Y137_SLICE_X23Y137_BQ),
.O(RIOB33_X105Y145_IOB_X1Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y147_OBUF (
.I(CLBLM_L_X16Y137_SLICE_X23Y137_CQ),
.O(RIOB33_X105Y147_IOB_X1Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y148_OBUF (
.I(CLBLM_L_X16Y139_SLICE_X22Y139_BQ),
.O(RIOB33_X105Y147_IOB_X1Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y149_IOB_X1Y149_OBUF (
.I(1'b1),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_OPAD)
  );
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A = CLBLL_L_X2Y116_SLICE_X0Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B = CLBLL_L_X2Y116_SLICE_X0Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C = CLBLL_L_X2Y116_SLICE_X0Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D = CLBLL_L_X2Y116_SLICE_X0Y116_DO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A = CLBLL_L_X2Y116_SLICE_X1Y116_AO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B = CLBLL_L_X2Y116_SLICE_X1Y116_BO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C = CLBLL_L_X2Y116_SLICE_X1Y116_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D = CLBLL_L_X2Y116_SLICE_X1Y116_DO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B = CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C = CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D = CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_AMUX = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A = CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B = CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C = CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D = CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A = CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B = CLBLL_L_X2Y132_SLICE_X0Y132_BO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C = CLBLL_L_X2Y132_SLICE_X0Y132_CO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D = CLBLL_L_X2Y132_SLICE_X0Y132_DO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A = CLBLL_L_X2Y132_SLICE_X1Y132_AO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B = CLBLL_L_X2Y132_SLICE_X1Y132_BO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C = CLBLL_L_X2Y132_SLICE_X1Y132_CO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D = CLBLL_L_X2Y132_SLICE_X1Y132_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C = CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D = CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A = CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B = CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C = CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D = CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A = CLBLL_L_X2Y135_SLICE_X0Y135_AO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B = CLBLL_L_X2Y135_SLICE_X0Y135_BO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C = CLBLL_L_X2Y135_SLICE_X0Y135_CO6;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D = CLBLL_L_X2Y135_SLICE_X0Y135_DO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A = CLBLL_L_X2Y135_SLICE_X1Y135_AO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B = CLBLL_L_X2Y135_SLICE_X1Y135_BO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C = CLBLL_L_X2Y135_SLICE_X1Y135_CO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D = CLBLL_L_X2Y135_SLICE_X1Y135_DO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_AMUX = CLBLL_L_X2Y135_SLICE_X1Y135_A5Q;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A = CLBLL_L_X2Y137_SLICE_X0Y137_AO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C = CLBLL_L_X2Y137_SLICE_X0Y137_CO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D = CLBLL_L_X2Y137_SLICE_X0Y137_DO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_AMUX = CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A = CLBLL_L_X2Y137_SLICE_X1Y137_AO6;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B = CLBLL_L_X2Y137_SLICE_X1Y137_BO6;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C = CLBLL_L_X2Y137_SLICE_X1Y137_CO6;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D = CLBLL_L_X2Y137_SLICE_X1Y137_DO6;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_AMUX = CLBLL_L_X2Y137_SLICE_X1Y137_AO5;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_BMUX = CLBLL_L_X2Y137_SLICE_X1Y137_BO5;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B = CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C = CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D = CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_AMUX = CLBLL_L_X2Y138_SLICE_X0Y138_A_XOR;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_BMUX = CLBLL_L_X2Y138_SLICE_X0Y138_B_XOR;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_CMUX = CLBLL_L_X2Y138_SLICE_X0Y138_C_XOR;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_DMUX = CLBLL_L_X2Y138_SLICE_X0Y138_D_XOR;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A = CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B = CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C = CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D = CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_AMUX = CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A = CLBLL_L_X2Y139_SLICE_X0Y139_AO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B = CLBLL_L_X2Y139_SLICE_X0Y139_BO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C = CLBLL_L_X2Y139_SLICE_X0Y139_CO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D = CLBLL_L_X2Y139_SLICE_X0Y139_DO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_AMUX = CLBLL_L_X2Y139_SLICE_X0Y139_A_XOR;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_BMUX = CLBLL_L_X2Y139_SLICE_X0Y139_B_XOR;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_CMUX = CLBLL_L_X2Y139_SLICE_X0Y139_C_XOR;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_DMUX = CLBLL_L_X2Y139_SLICE_X0Y139_D_XOR;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A = CLBLL_L_X2Y139_SLICE_X1Y139_AO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B = CLBLL_L_X2Y139_SLICE_X1Y139_BO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C = CLBLL_L_X2Y139_SLICE_X1Y139_CO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D = CLBLL_L_X2Y139_SLICE_X1Y139_DO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_AMUX = CLBLL_L_X2Y139_SLICE_X1Y139_AO5;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_BMUX = CLBLL_L_X2Y139_SLICE_X1Y139_BO5;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_CMUX = CLBLL_L_X2Y139_SLICE_X1Y139_CO5;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_DMUX = CLBLL_L_X2Y139_SLICE_X1Y139_DO5;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A = CLBLL_L_X2Y140_SLICE_X0Y140_AO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B = CLBLL_L_X2Y140_SLICE_X0Y140_BO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C = CLBLL_L_X2Y140_SLICE_X0Y140_CO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D = CLBLL_L_X2Y140_SLICE_X0Y140_DO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_AMUX = CLBLL_L_X2Y140_SLICE_X0Y140_A_XOR;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_BMUX = CLBLL_L_X2Y140_SLICE_X0Y140_B_XOR;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_CMUX = CLBLL_L_X2Y140_SLICE_X0Y140_C_XOR;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_DMUX = CLBLL_L_X2Y140_SLICE_X0Y140_D_XOR;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B = CLBLL_L_X2Y140_SLICE_X1Y140_BO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C = CLBLL_L_X2Y140_SLICE_X1Y140_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D = CLBLL_L_X2Y140_SLICE_X1Y140_DO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A = CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B = CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C = CLBLL_L_X2Y141_SLICE_X0Y141_CO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D = CLBLL_L_X2Y141_SLICE_X0Y141_DO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_AMUX = CLBLL_L_X2Y141_SLICE_X0Y141_A_XOR;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_BMUX = CLBLL_L_X2Y141_SLICE_X0Y141_B_XOR;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_CMUX = CLBLL_L_X2Y141_SLICE_X0Y141_C_XOR;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B = CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C = CLBLL_L_X2Y141_SLICE_X1Y141_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D = CLBLL_L_X2Y141_SLICE_X1Y141_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_DMUX = CLBLL_L_X2Y141_SLICE_X1Y141_D_XOR;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A = CLBLL_L_X2Y142_SLICE_X0Y142_AO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B = CLBLL_L_X2Y142_SLICE_X0Y142_BO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D = CLBLL_L_X2Y142_SLICE_X0Y142_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A = CLBLL_L_X2Y142_SLICE_X1Y142_AO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B = CLBLL_L_X2Y142_SLICE_X1Y142_BO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C = CLBLL_L_X2Y142_SLICE_X1Y142_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D = CLBLL_L_X2Y142_SLICE_X1Y142_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_CMUX = CLBLL_L_X2Y142_SLICE_X1Y142_C_XOR;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_DMUX = CLBLL_L_X2Y142_SLICE_X1Y142_D_XOR;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A = CLBLL_L_X2Y143_SLICE_X0Y143_AO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B = CLBLL_L_X2Y143_SLICE_X0Y143_BO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C = CLBLL_L_X2Y143_SLICE_X0Y143_CO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D = CLBLL_L_X2Y143_SLICE_X0Y143_DO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A = CLBLL_L_X2Y143_SLICE_X1Y143_AO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B = CLBLL_L_X2Y143_SLICE_X1Y143_BO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C = CLBLL_L_X2Y143_SLICE_X1Y143_CO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D = CLBLL_L_X2Y143_SLICE_X1Y143_DO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A = CLBLL_L_X2Y144_SLICE_X0Y144_AO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B = CLBLL_L_X2Y144_SLICE_X0Y144_BO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C = CLBLL_L_X2Y144_SLICE_X0Y144_CO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D = CLBLL_L_X2Y144_SLICE_X0Y144_DO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_AMUX = CLBLL_L_X2Y144_SLICE_X0Y144_A5Q;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A = CLBLL_L_X2Y144_SLICE_X1Y144_AO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B = CLBLL_L_X2Y144_SLICE_X1Y144_BO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C = CLBLL_L_X2Y144_SLICE_X1Y144_CO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D = CLBLL_L_X2Y144_SLICE_X1Y144_DO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_AMUX = CLBLL_L_X2Y144_SLICE_X1Y144_AO5;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A = CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B = CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C = CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D = CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_AMUX = CLBLL_L_X2Y145_SLICE_X0Y145_A5Q;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A = CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B = CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C = CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D = CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B = CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C = CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D = CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_AMUX = CLBLL_L_X2Y147_SLICE_X0Y147_A5Q;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C = CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D = CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A = CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B = CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C = CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D = CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D = CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_AMUX = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A = CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B = CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C = CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D = CLBLL_L_X2Y149_SLICE_X0Y149_DO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A = CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B = CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C = CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D = CLBLL_L_X2Y149_SLICE_X1Y149_DO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A = CLBLL_L_X2Y152_SLICE_X0Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B = CLBLL_L_X2Y152_SLICE_X0Y152_BO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C = CLBLL_L_X2Y152_SLICE_X0Y152_CO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D = CLBLL_L_X2Y152_SLICE_X0Y152_DO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C = CLBLL_L_X2Y152_SLICE_X1Y152_CO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D = CLBLL_L_X2Y152_SLICE_X1Y152_DO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A = CLBLL_L_X2Y153_SLICE_X0Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B = CLBLL_L_X2Y153_SLICE_X0Y153_BO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C = CLBLL_L_X2Y153_SLICE_X0Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D = CLBLL_L_X2Y153_SLICE_X0Y153_DO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_AMUX = CLBLL_L_X2Y153_SLICE_X0Y153_A5Q;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_BMUX = CLBLL_L_X2Y153_SLICE_X0Y153_B5Q;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_CMUX = CLBLL_L_X2Y153_SLICE_X0Y153_C5Q;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_DMUX = CLBLL_L_X2Y153_SLICE_X0Y153_D5Q;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A = CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_AMUX = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A = CLBLL_L_X2Y155_SLICE_X0Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B = CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C = CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D = CLBLL_L_X2Y155_SLICE_X0Y155_DO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A = CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_A = CLBLL_L_X2Y156_SLICE_X0Y156_AO6;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_B = CLBLL_L_X2Y156_SLICE_X0Y156_BO6;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_C = CLBLL_L_X2Y156_SLICE_X0Y156_CO6;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_D = CLBLL_L_X2Y156_SLICE_X0Y156_DO6;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_A = CLBLL_L_X2Y156_SLICE_X1Y156_AO6;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_B = CLBLL_L_X2Y156_SLICE_X1Y156_BO6;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_C = CLBLL_L_X2Y156_SLICE_X1Y156_CO6;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_D = CLBLL_L_X2Y156_SLICE_X1Y156_DO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A = CLBLL_L_X2Y157_SLICE_X0Y157_AO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B = CLBLL_L_X2Y157_SLICE_X0Y157_BO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C = CLBLL_L_X2Y157_SLICE_X0Y157_CO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D = CLBLL_L_X2Y157_SLICE_X0Y157_DO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_BMUX = CLBLL_L_X2Y157_SLICE_X0Y157_BO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A = CLBLL_L_X2Y157_SLICE_X1Y157_AO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B = CLBLL_L_X2Y157_SLICE_X1Y157_BO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C = CLBLL_L_X2Y157_SLICE_X1Y157_CO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D = CLBLL_L_X2Y157_SLICE_X1Y157_DO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A = CLBLL_L_X2Y158_SLICE_X0Y158_AO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B = CLBLL_L_X2Y158_SLICE_X0Y158_BO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C = CLBLL_L_X2Y158_SLICE_X0Y158_CO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D = CLBLL_L_X2Y158_SLICE_X0Y158_DO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_AMUX = CLBLL_L_X2Y158_SLICE_X0Y158_A5Q;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A = CLBLL_L_X2Y158_SLICE_X1Y158_AO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B = CLBLL_L_X2Y158_SLICE_X1Y158_BO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C = CLBLL_L_X2Y158_SLICE_X1Y158_CO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D = CLBLL_L_X2Y158_SLICE_X1Y158_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B = CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_AMUX = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B = CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B = CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C = CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A = CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A = CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_AMUX = CLBLL_L_X4Y133_SLICE_X5Y133_F7AMUX_O;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_DMUX = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B = CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_AMUX = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_AMUX = CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A = CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B = CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C = CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D = CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_AMUX = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_BMUX = CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_CMUX = CLBLL_L_X4Y135_SLICE_X4Y135_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_DMUX = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A = CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B = CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C = CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_AMUX = CLBLL_L_X4Y135_SLICE_X5Y135_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_BMUX = CLBLL_L_X4Y135_SLICE_X5Y135_B5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_CMUX = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_DMUX = CLBLL_L_X4Y135_SLICE_X5Y135_DO5;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A = CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B = CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C = CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D = CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A = CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D = CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_AMUX = CLBLL_L_X4Y136_SLICE_X5Y136_AO5;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_BMUX = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B = CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C = CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D = CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_AMUX = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A = CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B = CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C = CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D = CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_BMUX = CLBLL_L_X4Y137_SLICE_X5Y137_BO5;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A = CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B = CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C = CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_AMUX = CLBLL_L_X4Y138_SLICE_X5Y138_AO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_AMUX = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A = CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B = CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_AMUX = CLBLL_L_X4Y141_SLICE_X4Y141_F7AMUX_O;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_CMUX = CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_DMUX = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A = CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_BMUX = CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_CMUX = CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_DMUX = CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A = CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AMUX = CLBLL_L_X4Y142_SLICE_X4Y142_F7AMUX_O;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_CMUX = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_AMUX = CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_BMUX = CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CMUX = CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_DMUX = CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_AMUX = CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_BMUX = CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CMUX = CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_DMUX = CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C = CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_AMUX = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A = CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B = CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C = CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D = CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_AMUX = CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_BMUX = CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CMUX = CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_DMUX = CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_AMUX = CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_CMUX = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A = CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_AMUX = CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A = CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A = CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B = CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_AMUX = CLBLL_L_X4Y147_SLICE_X5Y147_AO5;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_AMUX = CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A = CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B = CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C = CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_AMUX = CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A = CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B = CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_AMUX = CLBLL_L_X4Y149_SLICE_X4Y149_AO5;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_CMUX = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_DMUX = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A = CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_AMUX = CLBLL_L_X4Y149_SLICE_X5Y149_AO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_BMUX = CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_CMUX = CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_AMUX = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A = CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B = CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C = CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D = CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_AMUX = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A = CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B = CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D = CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_DMUX = CLBLL_L_X4Y151_SLICE_X4Y151_DO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A = CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B = CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C = CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D = CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A = CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B = CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C = CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D = CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B = CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C = CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A = CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C = CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D = CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A = CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B = CLBLL_L_X4Y155_SLICE_X5Y155_BO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C = CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D = CLBLL_L_X4Y155_SLICE_X5Y155_DO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A = CLBLL_L_X4Y156_SLICE_X4Y156_AO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B = CLBLL_L_X4Y156_SLICE_X4Y156_BO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D = CLBLL_L_X4Y156_SLICE_X4Y156_DO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A = CLBLL_L_X4Y156_SLICE_X5Y156_AO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B = CLBLL_L_X4Y156_SLICE_X5Y156_BO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C = CLBLL_L_X4Y156_SLICE_X5Y156_CO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D = CLBLL_L_X4Y156_SLICE_X5Y156_DO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_A = CLBLL_L_X26Y133_SLICE_X38Y133_AO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_B = CLBLL_L_X26Y133_SLICE_X38Y133_BO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_C = CLBLL_L_X26Y133_SLICE_X38Y133_CO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_D = CLBLL_L_X26Y133_SLICE_X38Y133_DO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_AMUX = CLBLL_L_X26Y133_SLICE_X38Y133_AO5;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_BMUX = CLBLL_L_X26Y133_SLICE_X38Y133_BO5;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_CMUX = CLBLL_L_X26Y133_SLICE_X38Y133_CO5;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_DMUX = CLBLL_L_X26Y133_SLICE_X38Y133_DO5;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_A = CLBLL_L_X26Y133_SLICE_X39Y133_AO6;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_B = CLBLL_L_X26Y133_SLICE_X39Y133_BO6;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_C = CLBLL_L_X26Y133_SLICE_X39Y133_CO6;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_D = CLBLL_L_X26Y133_SLICE_X39Y133_DO6;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_A = CLBLL_L_X26Y135_SLICE_X38Y135_AO6;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_B = CLBLL_L_X26Y135_SLICE_X38Y135_BO6;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_C = CLBLL_L_X26Y135_SLICE_X38Y135_CO6;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_D = CLBLL_L_X26Y135_SLICE_X38Y135_DO6;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_AMUX = CLBLL_L_X26Y135_SLICE_X38Y135_AO5;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_A = CLBLL_L_X26Y135_SLICE_X39Y135_AO6;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_B = CLBLL_L_X26Y135_SLICE_X39Y135_BO6;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_C = CLBLL_L_X26Y135_SLICE_X39Y135_CO6;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_D = CLBLL_L_X26Y135_SLICE_X39Y135_DO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A = CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B = CLBLL_L_X26Y136_SLICE_X38Y136_BO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C = CLBLL_L_X26Y136_SLICE_X38Y136_CO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D = CLBLL_L_X26Y136_SLICE_X38Y136_DO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_AMUX = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_BMUX = CLBLL_L_X26Y136_SLICE_X38Y136_BO5;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A = CLBLL_L_X26Y136_SLICE_X39Y136_AO6;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B = CLBLL_L_X26Y136_SLICE_X39Y136_BO6;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C = CLBLL_L_X26Y136_SLICE_X39Y136_CO6;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D = CLBLL_L_X26Y136_SLICE_X39Y136_DO6;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_A = CLBLL_L_X26Y138_SLICE_X38Y138_AO6;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_B = CLBLL_L_X26Y138_SLICE_X38Y138_BO6;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_C = CLBLL_L_X26Y138_SLICE_X38Y138_CO6;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_D = CLBLL_L_X26Y138_SLICE_X38Y138_DO6;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_AMUX = CLBLL_L_X26Y138_SLICE_X38Y138_AO5;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_A = CLBLL_L_X26Y138_SLICE_X39Y138_AO6;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_B = CLBLL_L_X26Y138_SLICE_X39Y138_BO6;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_C = CLBLL_L_X26Y138_SLICE_X39Y138_CO6;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_D = CLBLL_L_X26Y138_SLICE_X39Y138_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_AMUX = CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_BMUX = CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A = CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_BMUX = CLBLM_L_X8Y134_SLICE_X10Y134_F8MUX_O;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B = CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A = CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A = CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A = CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_CMUX = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A = CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B = CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_BMUX = CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_CMUX = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A = CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B = CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D = CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_AMUX = CLBLM_L_X8Y137_SLICE_X10Y137_AO5;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_CMUX = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A = CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B = CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_CMUX = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C = CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_BMUX = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A = CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_AMUX = CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C = CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D = CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_AMUX = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A = CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B = CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_AMUX = CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A = CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B = CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_CMUX = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_DMUX = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_AMUX = CLBLM_L_X8Y140_SLICE_X11Y140_AO5;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_BMUX = CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_CMUX = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B = CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_AMUX = CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_BMUX = CLBLM_L_X8Y141_SLICE_X10Y141_BO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A = CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C = CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_AMUX = CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_DMUX = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A = CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_BMUX = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_AMUX = CLBLM_L_X8Y142_SLICE_X11Y142_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A = CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CMUX = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_DMUX = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_BMUX = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_BMUX = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_AMUX = CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A = CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B = CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_AMUX = CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A = CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B = CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C = CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_AMUX = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A = CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B = CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C = CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D = CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_CMUX = CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A = CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D = CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A = CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B = CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_AMUX = CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A = CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B = CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B = CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_AMUX = CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_CMUX = CLBLM_L_X8Y149_SLICE_X10Y149_CO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_DMUX = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A = CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B = CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C = CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_AMUX = CLBLM_L_X8Y149_SLICE_X11Y149_F7AMUX_O;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A = CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C = CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A = CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B = CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D = CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_BMUX = CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A = CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_AMUX = CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_BMUX = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_AMUX = CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_BMUX = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_DMUX = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_BMUX = CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CMUX = CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_AMUX = CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A = CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A = CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_AMUX = CLBLM_L_X10Y133_SLICE_X13Y133_AO5;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A = CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B = CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A = CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_AMUX = CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_BMUX = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B = CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_AMUX = CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_AMUX = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_BMUX = CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A = CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_BMUX = CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CMUX = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_AMUX = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_BMUX = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_AMUX = CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_AMUX = CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_BMUX = CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_CMUX = CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_DMUX = CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A = CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D = CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A = CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D = CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_AMUX = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A = CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C = CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D = CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A = CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B = CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_AMUX = CLBLM_L_X10Y140_SLICE_X12Y140_AO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A = CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B = CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C = CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A = CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C = CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A = CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B = CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_CMUX = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_AMUX = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A = CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_AMUX = CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_BMUX = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_BMUX = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_AMUX = CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_BMUX = CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_CMUX = CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_DMUX = CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_DMUX = CLBLM_L_X10Y144_SLICE_X13Y144_DO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_AMUX = CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_BMUX = CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CMUX = CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_DMUX = CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_DMUX = CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A = CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B = CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C = CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_AMUX = CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_BMUX = CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CMUX = CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_DMUX = CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A = CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_AMUX = CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_BMUX = CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CMUX = CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A = CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_AMUX = CLBLM_L_X10Y147_SLICE_X13Y147_AO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_DMUX = CLBLM_L_X10Y147_SLICE_X13Y147_DO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A = CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_AMUX = CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A = CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B = CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D = CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A = CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A = CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C = CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A = CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C = CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_AMUX = CLBLM_L_X10Y150_SLICE_X13Y150_AO5;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_AMUX = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A = CLBLM_L_X12Y128_SLICE_X16Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C = CLBLM_L_X12Y128_SLICE_X16Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D = CLBLM_L_X12Y128_SLICE_X16Y128_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_BMUX = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A = CLBLM_L_X12Y128_SLICE_X17Y128_AO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B = CLBLM_L_X12Y128_SLICE_X17Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C = CLBLM_L_X12Y128_SLICE_X17Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D = CLBLM_L_X12Y128_SLICE_X17Y128_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A = CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B = CLBLM_L_X12Y129_SLICE_X16Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D = CLBLM_L_X12Y129_SLICE_X16Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_AMUX = CLBLM_L_X12Y129_SLICE_X16Y129_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A = CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D = CLBLM_L_X12Y129_SLICE_X17Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_AMUX = CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A = CLBLM_L_X12Y130_SLICE_X16Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B = CLBLM_L_X12Y130_SLICE_X16Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C = CLBLM_L_X12Y130_SLICE_X16Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D = CLBLM_L_X12Y130_SLICE_X17Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_AMUX = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_AMUX = CLBLM_L_X12Y131_SLICE_X16Y131_A5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_BMUX = CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_CMUX = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A = CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D = CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_AMUX = CLBLM_L_X12Y131_SLICE_X17Y131_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C = CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_AMUX = CLBLM_L_X12Y132_SLICE_X16Y132_AO5;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_BMUX = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_CMUX = CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A = CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B = CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D = CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_AMUX = CLBLM_L_X12Y132_SLICE_X17Y132_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_BMUX = CLBLM_L_X12Y132_SLICE_X17Y132_B5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_CMUX = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A = CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B = CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C = CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_BMUX = CLBLM_L_X12Y133_SLICE_X16Y133_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_DMUX = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B = CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C = CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_BMUX = CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B = CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C = CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_AMUX = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_BMUX = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_CMUX = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C = CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D = CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_AMUX = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A = CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C = CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D = CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B = CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_AMUX = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_CMUX = CLBLM_L_X12Y137_SLICE_X16Y137_CO5;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A = CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B = CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C = CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_CMUX = CLBLM_L_X12Y137_SLICE_X17Y137_CO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A = CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C = CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D = CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A = CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C = CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B = CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C = CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D = CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B = CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C = CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_DMUX = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A = CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B = CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C = CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D = CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_CMUX = CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A = CLBLM_L_X12Y140_SLICE_X17Y140_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B = CLBLM_L_X12Y140_SLICE_X17Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C = CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_DMUX = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A = CLBLM_L_X12Y141_SLICE_X16Y141_AO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B = CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C = CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D = CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_CMUX = CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A = CLBLM_L_X12Y141_SLICE_X17Y141_AO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B = CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C = CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_AMUX = CLBLM_L_X12Y141_SLICE_X17Y141_AO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A = CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B = CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C = CLBLM_L_X12Y142_SLICE_X16Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D = CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A = CLBLM_L_X12Y142_SLICE_X17Y142_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B = CLBLM_L_X12Y142_SLICE_X17Y142_BO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C = CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_AMUX = CLBLM_L_X12Y142_SLICE_X17Y142_AO5;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_DMUX = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B = CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C = CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_BMUX = CLBLM_L_X12Y143_SLICE_X16Y143_BO5;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A = CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B = CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C = CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B = CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C = CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_AMUX = CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_BMUX = CLBLM_L_X12Y144_SLICE_X16Y144_BO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A = CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B = CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C = CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D = CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_AMUX = CLBLM_L_X12Y144_SLICE_X17Y144_F7AMUX_O;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_CMUX = CLBLM_L_X12Y144_SLICE_X17Y144_CO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C = CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_AMUX = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B = CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_CMUX = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_DMUX = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D = CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A = CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B = CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_AMUX = CLBLM_L_X12Y146_SLICE_X17Y146_F7AMUX_O;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_CMUX = CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A = CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B = CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C = CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_AMUX = CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_BMUX = CLBLM_L_X12Y147_SLICE_X16Y147_B_XOR;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_CMUX = CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_DMUX = CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B = CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C = CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_AMUX = CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_BMUX = CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_CMUX = CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_DMUX = CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C = CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D = CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_AMUX = CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_BMUX = CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_CMUX = CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_DMUX = CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A = CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B = CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C = CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D = CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_AMUX = CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_BMUX = CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_CMUX = CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_DMUX = CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A = CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B = CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_AMUX = CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_BMUX = CLBLM_L_X12Y149_SLICE_X16Y149_B_CY;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A = CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B = CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_AMUX = CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_BMUX = CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_CMUX = CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_DMUX = CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C = CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D = CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_AMUX = CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A = CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B = CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C = CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D = CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_AMUX = CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_BMUX = CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_CMUX = CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A = CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_DMUX = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B = CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C = CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_BMUX = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_A = CLBLM_L_X16Y131_SLICE_X22Y131_AO6;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_B = CLBLM_L_X16Y131_SLICE_X22Y131_BO6;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_C = CLBLM_L_X16Y131_SLICE_X22Y131_CO6;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_D = CLBLM_L_X16Y131_SLICE_X22Y131_DO6;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_A = CLBLM_L_X16Y131_SLICE_X23Y131_AO6;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_B = CLBLM_L_X16Y131_SLICE_X23Y131_BO6;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_C = CLBLM_L_X16Y131_SLICE_X23Y131_CO6;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_D = CLBLM_L_X16Y131_SLICE_X23Y131_DO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_A = CLBLM_L_X16Y133_SLICE_X22Y133_AO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_B = CLBLM_L_X16Y133_SLICE_X22Y133_BO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_C = CLBLM_L_X16Y133_SLICE_X22Y133_CO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_D = CLBLM_L_X16Y133_SLICE_X22Y133_DO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_A = CLBLM_L_X16Y133_SLICE_X23Y133_AO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_B = CLBLM_L_X16Y133_SLICE_X23Y133_BO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_C = CLBLM_L_X16Y133_SLICE_X23Y133_CO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_D = CLBLM_L_X16Y133_SLICE_X23Y133_DO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_A = CLBLM_L_X16Y134_SLICE_X22Y134_AO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_B = CLBLM_L_X16Y134_SLICE_X22Y134_BO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_C = CLBLM_L_X16Y134_SLICE_X22Y134_CO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_D = CLBLM_L_X16Y134_SLICE_X22Y134_DO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_AMUX = CLBLM_L_X16Y134_SLICE_X22Y134_AO5;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_A = CLBLM_L_X16Y134_SLICE_X23Y134_AO6;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_B = CLBLM_L_X16Y134_SLICE_X23Y134_BO6;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_C = CLBLM_L_X16Y134_SLICE_X23Y134_CO6;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_D = CLBLM_L_X16Y134_SLICE_X23Y134_DO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A = CLBLM_L_X16Y135_SLICE_X22Y135_AO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B = CLBLM_L_X16Y135_SLICE_X22Y135_BO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C = CLBLM_L_X16Y135_SLICE_X22Y135_CO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D = CLBLM_L_X16Y135_SLICE_X22Y135_DO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A = CLBLM_L_X16Y135_SLICE_X23Y135_AO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B = CLBLM_L_X16Y135_SLICE_X23Y135_BO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C = CLBLM_L_X16Y135_SLICE_X23Y135_CO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D = CLBLM_L_X16Y135_SLICE_X23Y135_DO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B = CLBLM_L_X16Y136_SLICE_X22Y136_BO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C = CLBLM_L_X16Y136_SLICE_X22Y136_CO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D = CLBLM_L_X16Y136_SLICE_X22Y136_DO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_AMUX = CLBLM_L_X16Y136_SLICE_X22Y136_AO5;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A = CLBLM_L_X16Y136_SLICE_X23Y136_AO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B = CLBLM_L_X16Y136_SLICE_X23Y136_BO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C = CLBLM_L_X16Y136_SLICE_X23Y136_CO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D = CLBLM_L_X16Y136_SLICE_X23Y136_DO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A = CLBLM_L_X16Y137_SLICE_X22Y137_AO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B = CLBLM_L_X16Y137_SLICE_X22Y137_BO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C = CLBLM_L_X16Y137_SLICE_X22Y137_CO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D = CLBLM_L_X16Y137_SLICE_X22Y137_DO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_AMUX = CLBLM_L_X16Y137_SLICE_X22Y137_AO5;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_BMUX = CLBLM_L_X16Y137_SLICE_X22Y137_BO5;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A = CLBLM_L_X16Y137_SLICE_X23Y137_AO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B = CLBLM_L_X16Y137_SLICE_X23Y137_BO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C = CLBLM_L_X16Y137_SLICE_X23Y137_CO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D = CLBLM_L_X16Y137_SLICE_X23Y137_DO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_AMUX = CLBLM_L_X16Y137_SLICE_X23Y137_AO5;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_A = CLBLM_L_X16Y138_SLICE_X22Y138_AO6;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_B = CLBLM_L_X16Y138_SLICE_X22Y138_BO6;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_C = CLBLM_L_X16Y138_SLICE_X22Y138_CO6;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_D = CLBLM_L_X16Y138_SLICE_X22Y138_DO6;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_A = CLBLM_L_X16Y138_SLICE_X23Y138_AO6;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_B = CLBLM_L_X16Y138_SLICE_X23Y138_BO6;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_C = CLBLM_L_X16Y138_SLICE_X23Y138_CO6;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_D = CLBLM_L_X16Y138_SLICE_X23Y138_DO6;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_A = CLBLM_L_X16Y139_SLICE_X22Y139_AO6;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_B = CLBLM_L_X16Y139_SLICE_X22Y139_BO6;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_C = CLBLM_L_X16Y139_SLICE_X22Y139_CO6;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_D = CLBLM_L_X16Y139_SLICE_X22Y139_DO6;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_A = CLBLM_L_X16Y139_SLICE_X23Y139_AO6;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_B = CLBLM_L_X16Y139_SLICE_X23Y139_BO6;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_C = CLBLM_L_X16Y139_SLICE_X23Y139_CO6;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_D = CLBLM_L_X16Y139_SLICE_X23Y139_DO6;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_A = CLBLM_L_X16Y140_SLICE_X22Y140_AO6;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_B = CLBLM_L_X16Y140_SLICE_X22Y140_BO6;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_C = CLBLM_L_X16Y140_SLICE_X22Y140_CO6;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_D = CLBLM_L_X16Y140_SLICE_X22Y140_DO6;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_A = CLBLM_L_X16Y140_SLICE_X23Y140_AO6;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_B = CLBLM_L_X16Y140_SLICE_X23Y140_BO6;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_C = CLBLM_L_X16Y140_SLICE_X23Y140_CO6;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_D = CLBLM_L_X16Y140_SLICE_X23Y140_DO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_A = CLBLM_L_X16Y141_SLICE_X22Y141_AO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_B = CLBLM_L_X16Y141_SLICE_X22Y141_BO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_C = CLBLM_L_X16Y141_SLICE_X22Y141_CO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_D = CLBLM_L_X16Y141_SLICE_X22Y141_DO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_AMUX = CLBLM_L_X16Y141_SLICE_X22Y141_AO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_BMUX = CLBLM_L_X16Y141_SLICE_X22Y141_BO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_A = CLBLM_L_X16Y141_SLICE_X23Y141_AO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_B = CLBLM_L_X16Y141_SLICE_X23Y141_BO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_C = CLBLM_L_X16Y141_SLICE_X23Y141_CO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_D = CLBLM_L_X16Y141_SLICE_X23Y141_DO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_A = CLBLM_L_X16Y142_SLICE_X22Y142_AO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_B = CLBLM_L_X16Y142_SLICE_X22Y142_BO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_C = CLBLM_L_X16Y142_SLICE_X22Y142_CO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_D = CLBLM_L_X16Y142_SLICE_X22Y142_DO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_AMUX = CLBLM_L_X16Y142_SLICE_X22Y142_AO5;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_A = CLBLM_L_X16Y142_SLICE_X23Y142_AO6;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_B = CLBLM_L_X16Y142_SLICE_X23Y142_BO6;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_C = CLBLM_L_X16Y142_SLICE_X23Y142_CO6;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_D = CLBLM_L_X16Y142_SLICE_X23Y142_DO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_A = CLBLM_L_X16Y143_SLICE_X22Y143_AO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_B = CLBLM_L_X16Y143_SLICE_X22Y143_BO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_C = CLBLM_L_X16Y143_SLICE_X22Y143_CO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_D = CLBLM_L_X16Y143_SLICE_X22Y143_DO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_AMUX = CLBLM_L_X16Y143_SLICE_X22Y143_AO6;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_A = CLBLM_L_X16Y143_SLICE_X23Y143_AO6;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_B = CLBLM_L_X16Y143_SLICE_X23Y143_BO6;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_C = CLBLM_L_X16Y143_SLICE_X23Y143_CO6;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_D = CLBLM_L_X16Y143_SLICE_X23Y143_DO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_A = CLBLM_L_X16Y150_SLICE_X22Y150_AO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_B = CLBLM_L_X16Y150_SLICE_X22Y150_BO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_C = CLBLM_L_X16Y150_SLICE_X22Y150_CO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_D = CLBLM_L_X16Y150_SLICE_X22Y150_DO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_AMUX = CLBLM_L_X16Y150_SLICE_X22Y150_A_XOR;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_BMUX = CLBLM_L_X16Y150_SLICE_X22Y150_B_XOR;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_CMUX = CLBLM_L_X16Y150_SLICE_X22Y150_C_XOR;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_DMUX = CLBLM_L_X16Y150_SLICE_X22Y150_D_XOR;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_A = CLBLM_L_X16Y150_SLICE_X23Y150_AO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_B = CLBLM_L_X16Y150_SLICE_X23Y150_BO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_C = CLBLM_L_X16Y150_SLICE_X23Y150_CO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_D = CLBLM_L_X16Y150_SLICE_X23Y150_DO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_AMUX = CLBLM_L_X16Y150_SLICE_X23Y150_AO5;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_BMUX = CLBLM_L_X16Y150_SLICE_X23Y150_BO5;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_CMUX = CLBLM_L_X16Y150_SLICE_X23Y150_CO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_DMUX = CLBLM_L_X16Y150_SLICE_X23Y150_DO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A = CLBLM_L_X16Y151_SLICE_X22Y151_AO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B = CLBLM_L_X16Y151_SLICE_X22Y151_BO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C = CLBLM_L_X16Y151_SLICE_X22Y151_CO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D = CLBLM_L_X16Y151_SLICE_X22Y151_DO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_AMUX = CLBLM_L_X16Y151_SLICE_X22Y151_A_XOR;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_BMUX = CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_CMUX = CLBLM_L_X16Y151_SLICE_X22Y151_C_XOR;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_DMUX = CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A = CLBLM_L_X16Y151_SLICE_X23Y151_AO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B = CLBLM_L_X16Y151_SLICE_X23Y151_BO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C = CLBLM_L_X16Y151_SLICE_X23Y151_CO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D = CLBLM_L_X16Y151_SLICE_X23Y151_DO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_CMUX = CLBLM_L_X16Y151_SLICE_X23Y151_CO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A = CLBLM_L_X16Y152_SLICE_X22Y152_AO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B = CLBLM_L_X16Y152_SLICE_X22Y152_BO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C = CLBLM_L_X16Y152_SLICE_X22Y152_CO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D = CLBLM_L_X16Y152_SLICE_X22Y152_DO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_AMUX = CLBLM_L_X16Y152_SLICE_X22Y152_A_XOR;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_BMUX = CLBLM_L_X16Y152_SLICE_X22Y152_B_XOR;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_CMUX = CLBLM_L_X16Y152_SLICE_X22Y152_C_XOR;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_DMUX = CLBLM_L_X16Y152_SLICE_X22Y152_D_XOR;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A = CLBLM_L_X16Y152_SLICE_X23Y152_AO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B = CLBLM_L_X16Y152_SLICE_X23Y152_BO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C = CLBLM_L_X16Y152_SLICE_X23Y152_CO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D = CLBLM_L_X16Y152_SLICE_X23Y152_DO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_DMUX = CLBLM_L_X16Y152_SLICE_X23Y152_DO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A = CLBLM_L_X16Y153_SLICE_X22Y153_AO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B = CLBLM_L_X16Y153_SLICE_X22Y153_BO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C = CLBLM_L_X16Y153_SLICE_X22Y153_CO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D = CLBLM_L_X16Y153_SLICE_X22Y153_DO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_AMUX = CLBLM_L_X16Y153_SLICE_X22Y153_A_XOR;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_BMUX = CLBLM_L_X16Y153_SLICE_X22Y153_B_XOR;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_CMUX = CLBLM_L_X16Y153_SLICE_X22Y153_C_XOR;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_DMUX = CLBLM_L_X16Y153_SLICE_X22Y153_D_XOR;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B = CLBLM_L_X16Y153_SLICE_X23Y153_BO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C = CLBLM_L_X16Y153_SLICE_X23Y153_CO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D = CLBLM_L_X16Y153_SLICE_X23Y153_DO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_AMUX = CLBLM_L_X16Y153_SLICE_X23Y153_AO5;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A = CLBLM_L_X16Y154_SLICE_X22Y154_AO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B = CLBLM_L_X16Y154_SLICE_X22Y154_BO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C = CLBLM_L_X16Y154_SLICE_X22Y154_CO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D = CLBLM_L_X16Y154_SLICE_X22Y154_DO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_AMUX = CLBLM_L_X16Y154_SLICE_X22Y154_A_CY;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A = CLBLM_L_X16Y154_SLICE_X23Y154_AO6;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B = CLBLM_L_X16Y154_SLICE_X23Y154_BO6;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C = CLBLM_L_X16Y154_SLICE_X23Y154_CO6;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D = CLBLM_L_X16Y154_SLICE_X23Y154_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_AMUX = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_AMUX = CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A = CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B = CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_DMUX = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A = CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B = CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D = CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A = CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B = CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D = CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_BMUX = CLBLM_R_X3Y133_SLICE_X2Y133_BO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_AMUX = CLBLM_R_X3Y133_SLICE_X3Y133_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_BMUX = CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_CMUX = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A = CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B = CLBLM_R_X3Y134_SLICE_X2Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C = CLBLM_R_X3Y134_SLICE_X2Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D = CLBLM_R_X3Y134_SLICE_X2Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A = CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B = CLBLM_R_X3Y134_SLICE_X3Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C = CLBLM_R_X3Y134_SLICE_X3Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_AMUX = CLBLM_R_X3Y134_SLICE_X3Y134_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_DMUX = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A = CLBLM_R_X3Y136_SLICE_X2Y136_AO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B = CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C = CLBLM_R_X3Y136_SLICE_X2Y136_CO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D = CLBLM_R_X3Y136_SLICE_X2Y136_DO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_AMUX = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A = CLBLM_R_X3Y136_SLICE_X3Y136_AO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B = CLBLM_R_X3Y136_SLICE_X3Y136_BO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C = CLBLM_R_X3Y136_SLICE_X3Y136_CO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D = CLBLM_R_X3Y136_SLICE_X3Y136_DO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A = CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B = CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C = CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D = CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_AMUX = CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A = CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B = CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C = CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D = CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A = CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B = CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C = CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D = CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A = CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B = CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C = CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D = CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A = CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B = CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C = CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D = CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A = CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C = CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D = CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A = CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B = CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C = CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_AMUX = CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_BMUX = CLBLM_R_X3Y140_SLICE_X2Y140_BO5;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_DMUX = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A = CLBLM_R_X3Y140_SLICE_X3Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B = CLBLM_R_X3Y140_SLICE_X3Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C = CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D = CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D = CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_AMUX = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_AMUX = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_CMUX = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_DMUX = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D = CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A = CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A = CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C = CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B = CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C = CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_AMUX = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_DMUX = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A = CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_AMUX = CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_BMUX = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A = CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B = CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C = CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D = CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C = CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D = CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_AMUX = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_BMUX = CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B = CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B = CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C = CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A = CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C = CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_BMUX = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_CMUX = CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B = CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_AMUX = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_BMUX = CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_AMUX = CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_BMUX = CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B = CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_DMUX = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C = CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_AMUX = CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_DMUX = CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_AMUX = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_BMUX = CLBLM_R_X3Y152_SLICE_X2Y152_BO5;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D = CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_AMUX = CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_BMUX = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_AMUX = CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B = CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C = CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D = CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B = CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C = CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D = CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A = CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_AMUX = CLBLM_R_X3Y155_SLICE_X2Y155_A5Q;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_CMUX = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_DMUX = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B = CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B = CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_AMUX = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A = CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B = CLBLM_R_X3Y156_SLICE_X3Y156_BO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C = CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D = CLBLM_R_X3Y156_SLICE_X3Y156_DO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A = CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B = CLBLM_R_X3Y157_SLICE_X2Y157_BO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C = CLBLM_R_X3Y157_SLICE_X2Y157_CO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D = CLBLM_R_X3Y157_SLICE_X2Y157_DO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A = CLBLM_R_X3Y157_SLICE_X3Y157_AO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B = CLBLM_R_X3Y157_SLICE_X3Y157_BO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C = CLBLM_R_X3Y157_SLICE_X3Y157_CO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D = CLBLM_R_X3Y157_SLICE_X3Y157_DO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B = CLBLM_R_X3Y158_SLICE_X2Y158_BO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C = CLBLM_R_X3Y158_SLICE_X2Y158_CO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D = CLBLM_R_X3Y158_SLICE_X2Y158_DO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_AMUX = CLBLM_R_X3Y158_SLICE_X2Y158_A5Q;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A = CLBLM_R_X3Y158_SLICE_X3Y158_AO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B = CLBLM_R_X3Y158_SLICE_X3Y158_BO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C = CLBLM_R_X3Y158_SLICE_X3Y158_CO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D = CLBLM_R_X3Y158_SLICE_X3Y158_DO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_BMUX = CLBLM_R_X3Y158_SLICE_X3Y158_BO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_CMUX = CLBLM_R_X3Y158_SLICE_X3Y158_CO6;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_A = CLBLM_R_X3Y159_SLICE_X2Y159_AO6;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_B = CLBLM_R_X3Y159_SLICE_X2Y159_BO6;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_C = CLBLM_R_X3Y159_SLICE_X2Y159_CO6;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_D = CLBLM_R_X3Y159_SLICE_X2Y159_DO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_A = CLBLM_R_X3Y159_SLICE_X3Y159_AO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_B = CLBLM_R_X3Y159_SLICE_X3Y159_BO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_C = CLBLM_R_X3Y159_SLICE_X3Y159_CO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_D = CLBLM_R_X3Y159_SLICE_X3Y159_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A = CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B = CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A = CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B = CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C = CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_AMUX = CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_BMUX = CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_CMUX = CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_DMUX = CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A = CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_AMUX = CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_BMUX = CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_CMUX = CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_DMUX = CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_BMUX = CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CMUX = CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_DMUX = CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_AMUX = CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_BMUX = CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CMUX = CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_DMUX = CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A = CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B = CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_AMUX = CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_BMUX = CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CMUX = CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_DMUX = CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A = CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B = CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C = CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_AMUX = CLBLM_R_X5Y131_SLICE_X7Y131_A_CY;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B = CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_AMUX = CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_BMUX = CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CMUX = CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_DMUX = CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A = CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A = CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_AMUX = CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_BMUX = CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_CMUX = CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_DMUX = CLBLM_R_X5Y133_SLICE_X6Y133_D_CY;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_AMUX = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_BMUX = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A = CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B = CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_CMUX = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A = CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_BMUX = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A = CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B = CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_DMUX = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B = CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C = CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_AMUX = CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B = CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_AMUX = CLBLM_R_X5Y137_SLICE_X6Y137_AO5;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A = CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B = CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C = CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_AMUX = CLBLM_R_X5Y137_SLICE_X7Y137_AO5;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_BMUX = CLBLM_R_X5Y137_SLICE_X7Y137_BO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C = CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_AMUX = CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A = CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B = CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_AMUX = CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_BMUX = CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_CMUX = CLBLM_R_X5Y138_SLICE_X7Y138_CO5;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A = CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A = CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B = CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_AMUX = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A = CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B = CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C = CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A = CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B = CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C = CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_AMUX = CLBLM_R_X5Y141_SLICE_X6Y141_F7AMUX_O;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B = CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_AMUX = CLBLM_R_X5Y141_SLICE_X7Y141_F7AMUX_O;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A = CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B = CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_AMUX = CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_BMUX = CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_CMUX = CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_DMUX = CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_AMUX = CLBLM_R_X5Y142_SLICE_X7Y142_F7AMUX_O;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CMUX = CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_DMUX = CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D = CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_AMUX = CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_BMUX = CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CMUX = CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_DMUX = CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_AMUX = CLBLM_R_X5Y143_SLICE_X7Y143_F7AMUX_O;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A = CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_AMUX = CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A = CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C = CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_AMUX = CLBLM_R_X5Y144_SLICE_X7Y144_AO5;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A = CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B = CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C = CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A = CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C = CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_AMUX = CLBLM_R_X5Y145_SLICE_X7Y145_AO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B = CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_AMUX = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A = CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B = CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C = CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B = CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_BMUX = CLBLM_R_X5Y147_SLICE_X6Y147_BO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_DMUX = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A = CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B = CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CMUX = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_AMUX = CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A = CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B = CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_AMUX = CLBLM_R_X5Y148_SLICE_X7Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_BMUX = CLBLM_R_X5Y148_SLICE_X7Y148_BO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_DMUX = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A = CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B = CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_AMUX = CLBLM_R_X5Y149_SLICE_X6Y149_AO5;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_CMUX = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A = CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B = CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C = CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B = CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D = CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A = CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_BMUX = CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_CMUX = CLBLM_R_X5Y150_SLICE_X7Y150_CO5;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_DMUX = CLBLM_R_X5Y150_SLICE_X7Y150_DO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B = CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C = CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D = CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_AMUX = CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_BMUX = CLBLM_R_X5Y151_SLICE_X6Y151_BO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_CMUX = CLBLM_R_X5Y151_SLICE_X6Y151_CO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A = CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_AMUX = CLBLM_R_X5Y151_SLICE_X7Y151_AO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_CMUX = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A = CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A = CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A = CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_BMUX = CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A = CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CMUX = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A = CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_BMUX = CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B = CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C = CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_AMUX = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A = CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C = CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A = CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B = CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C = CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_AMUX = CLBLM_R_X7Y134_SLICE_X8Y134_AO5;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A = CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B = CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_AMUX = CLBLM_R_X7Y134_SLICE_X9Y134_AO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_AMUX = CLBLM_R_X7Y135_SLICE_X8Y135_AO5;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A = CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B = CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_CMUX = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A = CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B = CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_BMUX = CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A = CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_AMUX = CLBLM_R_X7Y136_SLICE_X9Y136_AO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_BMUX = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B = CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_AMUX = CLBLM_R_X7Y137_SLICE_X8Y137_F7AMUX_O;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_CMUX = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_DMUX = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A = CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B = CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C = CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D = CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_AMUX = CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_BMUX = CLBLM_R_X7Y138_SLICE_X8Y138_B_XOR;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_CMUX = CLBLM_R_X7Y138_SLICE_X8Y138_C_XOR;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_DMUX = CLBLM_R_X7Y138_SLICE_X8Y138_D_XOR;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A = CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_AMUX = CLBLM_R_X7Y138_SLICE_X9Y138_AO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_AMUX = CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_BMUX = CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CMUX = CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_DMUX = CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A = CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_AMUX = CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_BMUX = CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A = CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B = CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C = CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_AMUX = CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_DMUX = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A = CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B = CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C = CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_AMUX = CLBLM_R_X7Y140_SLICE_X9Y140_F7AMUX_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A = CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_AMUX = CLBLM_R_X7Y141_SLICE_X8Y141_F7AMUX_O;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C = CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_AMUX = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_AMUX = CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A = CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C = CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_AMUX = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A = CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A = CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A = CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C = CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_AMUX = CLBLM_R_X7Y145_SLICE_X8Y145_AO5;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_BMUX = CLBLM_R_X7Y145_SLICE_X8Y145_BO5;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C = CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_AMUX = CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A = CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A = CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A = CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B = CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C = CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_BMUX = CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_AMUX = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_BMUX = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_CMUX = CLBLM_R_X7Y148_SLICE_X8Y148_CO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A = CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B = CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C = CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_AMUX = CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_DMUX = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A = CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B = CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C = CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D = CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_BMUX = CLBLM_R_X7Y149_SLICE_X8Y149_BO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A = CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_BMUX = CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A = CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B = CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A = CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_BMUX = CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B = CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C = CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_BMUX = CLBLM_R_X7Y151_SLICE_X8Y151_BO5;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A = CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B = CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C = CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C = CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_AMUX = CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_BMUX = CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_CMUX = CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_DMUX = CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A = CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_BMUX = CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_CMUX = CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_DMUX = CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_AMUX = CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_BMUX = CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CMUX = CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_DMUX = CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_AMUX = CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_BMUX = CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CMUX = CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_DMUX = CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A = CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_AMUX = CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_BMUX = CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CMUX = CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_DMUX = CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_AMUX = CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_BMUX = CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_CMUX = CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_DMUX = CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_AMUX = CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_BMUX = CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CMUX = CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_DMUX = CLBLM_R_X11Y133_SLICE_X14Y133_D_CY;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D = CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_AMUX = CLBLM_R_X11Y133_SLICE_X15Y133_A_CY;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CMUX = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D = CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C = CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_AMUX = CLBLM_R_X11Y135_SLICE_X15Y135_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B = CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_CMUX = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_BMUX = CLBLM_R_X11Y137_SLICE_X14Y137_F8MUX_O;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C = CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_AMUX = CLBLM_R_X11Y137_SLICE_X15Y137_AO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A = CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B = CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C = CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D = CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A = CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A = CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B = CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CMUX = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B = CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D = CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CMUX = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A = CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B = CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C = CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D = CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A = CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B = CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A = CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B = CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C = CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_AMUX = CLBLM_R_X11Y141_SLICE_X15Y141_AO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_BMUX = CLBLM_R_X11Y141_SLICE_X15Y141_BO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_CMUX = CLBLM_R_X11Y141_SLICE_X15Y141_CO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A = CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A = CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B = CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C = CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D = CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_AMUX = CLBLM_R_X11Y142_SLICE_X15Y142_F7AMUX_O;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_BMUX = CLBLM_R_X11Y142_SLICE_X15Y142_F8MUX_O;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_CMUX = CLBLM_R_X11Y142_SLICE_X15Y142_F7BMUX_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_BMUX = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A = CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_AMUX = CLBLM_R_X11Y143_SLICE_X15Y143_A5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_AMUX = CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_AMUX = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B = CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A = CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D = CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A = CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_DMUX = CLBLM_R_X11Y147_SLICE_X14Y147_DO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A = CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_AMUX = CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_BMUX = CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_CMUX = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_AMUX = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_AMUX = CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_BMUX = CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_AMUX = CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_AMUX = CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_BMUX = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A = CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B = CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_AMUX = CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A = CLBLM_R_X13Y128_SLICE_X18Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B = CLBLM_R_X13Y128_SLICE_X18Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D = CLBLM_R_X13Y128_SLICE_X18Y128_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_AMUX = CLBLM_R_X13Y128_SLICE_X18Y128_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_BMUX = CLBLM_R_X13Y128_SLICE_X18Y128_B5Q;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A = CLBLM_R_X13Y128_SLICE_X19Y128_AO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B = CLBLM_R_X13Y128_SLICE_X19Y128_BO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C = CLBLM_R_X13Y128_SLICE_X19Y128_CO6;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D = CLBLM_R_X13Y128_SLICE_X19Y128_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A = CLBLM_R_X13Y129_SLICE_X18Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B = CLBLM_R_X13Y129_SLICE_X18Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C = CLBLM_R_X13Y129_SLICE_X18Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_BMUX = CLBLM_R_X13Y129_SLICE_X18Y129_B5Q;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A = CLBLM_R_X13Y129_SLICE_X19Y129_AO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B = CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_BMUX = CLBLM_R_X13Y129_SLICE_X19Y129_BO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A = CLBLM_R_X13Y130_SLICE_X18Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B = CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A = CLBLM_R_X13Y130_SLICE_X19Y130_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D = CLBLM_R_X13Y130_SLICE_X19Y130_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A = CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B = CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C = CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D = CLBLM_R_X13Y131_SLICE_X18Y131_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_CMUX = CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A = CLBLM_R_X13Y131_SLICE_X19Y131_AO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B = CLBLM_R_X13Y131_SLICE_X19Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C = CLBLM_R_X13Y131_SLICE_X19Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D = CLBLM_R_X13Y131_SLICE_X19Y131_DO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C = CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D = CLBLM_R_X13Y132_SLICE_X18Y132_DO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_AMUX = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_BMUX = CLBLM_R_X13Y132_SLICE_X18Y132_BO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_CMUX = CLBLM_R_X13Y132_SLICE_X18Y132_CO5;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_DMUX = CLBLM_R_X13Y132_SLICE_X18Y132_D5Q;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A = CLBLM_R_X13Y132_SLICE_X19Y132_AO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B = CLBLM_R_X13Y132_SLICE_X19Y132_BO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C = CLBLM_R_X13Y132_SLICE_X19Y132_CO6;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D = CLBLM_R_X13Y132_SLICE_X19Y132_DO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A = CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B = CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C = CLBLM_R_X13Y133_SLICE_X18Y133_CO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D = CLBLM_R_X13Y133_SLICE_X18Y133_DO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_AMUX = CLBLM_R_X13Y133_SLICE_X18Y133_AO5;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_BMUX = CLBLM_R_X13Y133_SLICE_X18Y133_BO5;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A = CLBLM_R_X13Y133_SLICE_X19Y133_AO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B = CLBLM_R_X13Y133_SLICE_X19Y133_BO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D = CLBLM_R_X13Y133_SLICE_X19Y133_DO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_AMUX = CLBLM_R_X13Y133_SLICE_X19Y133_A5Q;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_BMUX = CLBLM_R_X13Y133_SLICE_X19Y133_B5Q;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_CMUX = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B = CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_AMUX = CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_BMUX = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_DMUX = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A = CLBLM_R_X13Y134_SLICE_X19Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B = CLBLM_R_X13Y134_SLICE_X19Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C = CLBLM_R_X13Y134_SLICE_X19Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D = CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_AMUX = CLBLM_R_X13Y134_SLICE_X19Y134_A5Q;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_BMUX = CLBLM_R_X13Y134_SLICE_X19Y134_B5Q;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_DMUX = CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A = CLBLM_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B = CLBLM_R_X13Y135_SLICE_X18Y135_BO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C = CLBLM_R_X13Y135_SLICE_X18Y135_CO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D = CLBLM_R_X13Y135_SLICE_X18Y135_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_AMUX = CLBLM_R_X13Y135_SLICE_X18Y135_AO5;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A = CLBLM_R_X13Y135_SLICE_X19Y135_AO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B = CLBLM_R_X13Y135_SLICE_X19Y135_BO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C = CLBLM_R_X13Y135_SLICE_X19Y135_CO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D = CLBLM_R_X13Y135_SLICE_X19Y135_DO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A = CLBLM_R_X13Y136_SLICE_X18Y136_AO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B = CLBLM_R_X13Y136_SLICE_X18Y136_BO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C = CLBLM_R_X13Y136_SLICE_X18Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D = CLBLM_R_X13Y136_SLICE_X18Y136_DO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_AMUX = CLBLM_R_X13Y136_SLICE_X18Y136_A5Q;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_BMUX = CLBLM_R_X13Y136_SLICE_X18Y136_B5Q;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A = CLBLM_R_X13Y136_SLICE_X19Y136_AO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B = CLBLM_R_X13Y136_SLICE_X19Y136_BO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C = CLBLM_R_X13Y136_SLICE_X19Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D = CLBLM_R_X13Y136_SLICE_X19Y136_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A = CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B = CLBLM_R_X13Y137_SLICE_X18Y137_BO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C = CLBLM_R_X13Y137_SLICE_X18Y137_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D = CLBLM_R_X13Y137_SLICE_X18Y137_DO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A = CLBLM_R_X13Y137_SLICE_X19Y137_AO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B = CLBLM_R_X13Y137_SLICE_X19Y137_BO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C = CLBLM_R_X13Y137_SLICE_X19Y137_CO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D = CLBLM_R_X13Y137_SLICE_X19Y137_DO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_AMUX = CLBLM_R_X13Y137_SLICE_X19Y137_AO5;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A = CLBLM_R_X13Y138_SLICE_X18Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C = CLBLM_R_X13Y138_SLICE_X18Y138_CO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D = CLBLM_R_X13Y138_SLICE_X18Y138_DO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_AMUX = CLBLM_R_X13Y138_SLICE_X18Y138_A5Q;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A = CLBLM_R_X13Y138_SLICE_X19Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B = CLBLM_R_X13Y138_SLICE_X19Y138_BO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C = CLBLM_R_X13Y138_SLICE_X19Y138_CO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A = CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C = CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D = CLBLM_R_X13Y139_SLICE_X18Y139_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C = CLBLM_R_X13Y139_SLICE_X19Y139_CO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_AMUX = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A = CLBLM_R_X13Y140_SLICE_X18Y140_AO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B = CLBLM_R_X13Y140_SLICE_X18Y140_BO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C = CLBLM_R_X13Y140_SLICE_X18Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D = CLBLM_R_X13Y140_SLICE_X18Y140_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_BMUX = CLBLM_R_X13Y140_SLICE_X18Y140_BO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A = CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B = CLBLM_R_X13Y140_SLICE_X19Y140_BO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C = CLBLM_R_X13Y140_SLICE_X19Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D = CLBLM_R_X13Y140_SLICE_X19Y140_DO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_AMUX = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_BMUX = CLBLM_R_X13Y140_SLICE_X19Y140_BO5;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A = CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D = CLBLM_R_X13Y141_SLICE_X18Y141_DO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_BMUX = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A = CLBLM_R_X13Y141_SLICE_X19Y141_AO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B = CLBLM_R_X13Y141_SLICE_X19Y141_BO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C = CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D = CLBLM_R_X13Y141_SLICE_X19Y141_DO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A = CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B = CLBLM_R_X13Y142_SLICE_X18Y142_BO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C = CLBLM_R_X13Y142_SLICE_X18Y142_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D = CLBLM_R_X13Y142_SLICE_X18Y142_DO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A = CLBLM_R_X13Y142_SLICE_X19Y142_AO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B = CLBLM_R_X13Y142_SLICE_X19Y142_BO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C = CLBLM_R_X13Y142_SLICE_X19Y142_CO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D = CLBLM_R_X13Y142_SLICE_X19Y142_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B = CLBLM_R_X13Y144_SLICE_X18Y144_BO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D = CLBLM_R_X13Y144_SLICE_X18Y144_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_AMUX = CLBLM_R_X13Y144_SLICE_X18Y144_A_XOR;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_BMUX = CLBLM_R_X13Y144_SLICE_X18Y144_B_XOR;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_CMUX = CLBLM_R_X13Y144_SLICE_X18Y144_C_XOR;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_DMUX = CLBLM_R_X13Y144_SLICE_X18Y144_D_XOR;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A = CLBLM_R_X13Y144_SLICE_X19Y144_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B = CLBLM_R_X13Y144_SLICE_X19Y144_BO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C = CLBLM_R_X13Y144_SLICE_X19Y144_CO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D = CLBLM_R_X13Y144_SLICE_X19Y144_DO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_AMUX = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_CMUX = CLBLM_R_X13Y144_SLICE_X19Y144_CO5;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A = CLBLM_R_X13Y145_SLICE_X18Y145_AO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B = CLBLM_R_X13Y145_SLICE_X18Y145_BO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C = CLBLM_R_X13Y145_SLICE_X18Y145_CO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D = CLBLM_R_X13Y145_SLICE_X18Y145_DO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_AMUX = CLBLM_R_X13Y145_SLICE_X18Y145_A_XOR;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_BMUX = CLBLM_R_X13Y145_SLICE_X18Y145_B_XOR;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_CMUX = CLBLM_R_X13Y145_SLICE_X18Y145_C_XOR;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_DMUX = CLBLM_R_X13Y145_SLICE_X18Y145_D_XOR;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A = CLBLM_R_X13Y145_SLICE_X19Y145_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B = CLBLM_R_X13Y145_SLICE_X19Y145_BO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D = CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_AMUX = CLBLM_R_X13Y145_SLICE_X19Y145_AO5;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_BMUX = CLBLM_R_X13Y145_SLICE_X19Y145_BO5;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A = CLBLM_R_X13Y146_SLICE_X18Y146_AO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B = CLBLM_R_X13Y146_SLICE_X18Y146_BO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C = CLBLM_R_X13Y146_SLICE_X18Y146_CO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D = CLBLM_R_X13Y146_SLICE_X18Y146_DO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_AMUX = CLBLM_R_X13Y146_SLICE_X18Y146_A_XOR;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_BMUX = CLBLM_R_X13Y146_SLICE_X18Y146_B_XOR;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_CMUX = CLBLM_R_X13Y146_SLICE_X18Y146_C_XOR;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_DMUX = CLBLM_R_X13Y146_SLICE_X18Y146_D_XOR;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B = CLBLM_R_X13Y146_SLICE_X19Y146_BO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C = CLBLM_R_X13Y146_SLICE_X19Y146_CO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D = CLBLM_R_X13Y146_SLICE_X19Y146_DO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_AMUX = CLBLM_R_X13Y146_SLICE_X19Y146_AO5;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A = CLBLM_R_X13Y147_SLICE_X18Y147_AO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B = CLBLM_R_X13Y147_SLICE_X18Y147_BO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C = CLBLM_R_X13Y147_SLICE_X18Y147_CO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D = CLBLM_R_X13Y147_SLICE_X18Y147_DO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_AMUX = CLBLM_R_X13Y147_SLICE_X18Y147_A_XOR;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_BMUX = CLBLM_R_X13Y147_SLICE_X18Y147_B_XOR;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_CMUX = CLBLM_R_X13Y147_SLICE_X18Y147_C_XOR;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A = CLBLM_R_X13Y147_SLICE_X19Y147_AO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C = CLBLM_R_X13Y147_SLICE_X19Y147_CO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D = CLBLM_R_X13Y147_SLICE_X19Y147_DO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_AMUX = CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_CMUX = CLBLM_R_X13Y147_SLICE_X19Y147_CO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_DMUX = CLBLM_R_X13Y147_SLICE_X19Y147_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A = CLBLM_R_X13Y148_SLICE_X18Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B = CLBLM_R_X13Y148_SLICE_X18Y148_BO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C = CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D = CLBLM_R_X13Y148_SLICE_X18Y148_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_AMUX = CLBLM_R_X13Y148_SLICE_X18Y148_AO5;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A = CLBLM_R_X13Y148_SLICE_X19Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B = CLBLM_R_X13Y148_SLICE_X19Y148_BO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C = CLBLM_R_X13Y148_SLICE_X19Y148_CO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D = CLBLM_R_X13Y148_SLICE_X19Y148_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B = CLBLM_R_X13Y149_SLICE_X18Y149_BO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C = CLBLM_R_X13Y149_SLICE_X18Y149_CO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D = CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_AMUX = CLBLM_R_X13Y149_SLICE_X18Y149_F7AMUX_O;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A = CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B = CLBLM_R_X13Y149_SLICE_X19Y149_BO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C = CLBLM_R_X13Y149_SLICE_X19Y149_CO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D = CLBLM_R_X13Y149_SLICE_X19Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_AMUX = CLBLM_R_X13Y149_SLICE_X19Y149_AO5;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B = CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C = CLBLM_R_X13Y150_SLICE_X18Y150_CO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D = CLBLM_R_X13Y150_SLICE_X18Y150_DO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A = CLBLM_R_X13Y150_SLICE_X19Y150_AO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B = CLBLM_R_X13Y150_SLICE_X19Y150_BO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C = CLBLM_R_X13Y150_SLICE_X19Y150_CO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D = CLBLM_R_X13Y150_SLICE_X19Y150_DO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_AMUX = CLBLM_R_X13Y150_SLICE_X19Y150_F7AMUX_O;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A = CLBLM_R_X15Y128_SLICE_X20Y128_AO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B = CLBLM_R_X15Y128_SLICE_X20Y128_BO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C = CLBLM_R_X15Y128_SLICE_X20Y128_CO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D = CLBLM_R_X15Y128_SLICE_X20Y128_DO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_AMUX = CLBLM_R_X15Y128_SLICE_X20Y128_A5Q;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_BMUX = CLBLM_R_X15Y128_SLICE_X20Y128_B5Q;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A = CLBLM_R_X15Y128_SLICE_X21Y128_AO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B = CLBLM_R_X15Y128_SLICE_X21Y128_BO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C = CLBLM_R_X15Y128_SLICE_X21Y128_CO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D = CLBLM_R_X15Y128_SLICE_X21Y128_DO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A = CLBLM_R_X15Y129_SLICE_X20Y129_AO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B = CLBLM_R_X15Y129_SLICE_X20Y129_BO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C = CLBLM_R_X15Y129_SLICE_X20Y129_CO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D = CLBLM_R_X15Y129_SLICE_X20Y129_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A = CLBLM_R_X15Y129_SLICE_X21Y129_AO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B = CLBLM_R_X15Y129_SLICE_X21Y129_BO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C = CLBLM_R_X15Y129_SLICE_X21Y129_CO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_BMUX = CLBLM_R_X15Y129_SLICE_X21Y129_B5Q;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A = CLBLM_R_X15Y130_SLICE_X20Y130_AO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B = CLBLM_R_X15Y130_SLICE_X20Y130_BO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C = CLBLM_R_X15Y130_SLICE_X20Y130_CO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D = CLBLM_R_X15Y130_SLICE_X20Y130_DO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_AMUX = CLBLM_R_X15Y130_SLICE_X20Y130_AO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A = CLBLM_R_X15Y130_SLICE_X21Y130_AO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B = CLBLM_R_X15Y130_SLICE_X21Y130_BO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C = CLBLM_R_X15Y130_SLICE_X21Y130_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D = CLBLM_R_X15Y130_SLICE_X21Y130_DO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A = CLBLM_R_X15Y131_SLICE_X20Y131_AO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B = CLBLM_R_X15Y131_SLICE_X20Y131_BO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C = CLBLM_R_X15Y131_SLICE_X20Y131_CO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D = CLBLM_R_X15Y131_SLICE_X20Y131_DO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A = CLBLM_R_X15Y131_SLICE_X21Y131_AO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B = CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C = CLBLM_R_X15Y131_SLICE_X21Y131_CO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D = CLBLM_R_X15Y131_SLICE_X21Y131_DO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_AMUX = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_BMUX = CLBLM_R_X15Y131_SLICE_X21Y131_BO5;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_A = CLBLM_R_X15Y133_SLICE_X20Y133_AO6;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_B = CLBLM_R_X15Y133_SLICE_X20Y133_BO6;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_C = CLBLM_R_X15Y133_SLICE_X20Y133_CO6;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_D = CLBLM_R_X15Y133_SLICE_X20Y133_DO6;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_A = CLBLM_R_X15Y133_SLICE_X21Y133_AO6;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_B = CLBLM_R_X15Y133_SLICE_X21Y133_BO6;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_C = CLBLM_R_X15Y133_SLICE_X21Y133_CO6;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_D = CLBLM_R_X15Y133_SLICE_X21Y133_DO6;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_A = CLBLM_R_X15Y134_SLICE_X20Y134_AO6;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_B = CLBLM_R_X15Y134_SLICE_X20Y134_BO6;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_C = CLBLM_R_X15Y134_SLICE_X20Y134_CO6;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_D = CLBLM_R_X15Y134_SLICE_X20Y134_DO6;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_AMUX = CLBLM_R_X15Y134_SLICE_X20Y134_A_XOR;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_BMUX = CLBLM_R_X15Y134_SLICE_X20Y134_B_XOR;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_CMUX = CLBLM_R_X15Y134_SLICE_X20Y134_C_XOR;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_DMUX = CLBLM_R_X15Y134_SLICE_X20Y134_D_XOR;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_A = CLBLM_R_X15Y134_SLICE_X21Y134_AO6;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_B = CLBLM_R_X15Y134_SLICE_X21Y134_BO6;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_C = CLBLM_R_X15Y134_SLICE_X21Y134_CO6;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_D = CLBLM_R_X15Y134_SLICE_X21Y134_DO6;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A = CLBLM_R_X15Y135_SLICE_X20Y135_AO6;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B = CLBLM_R_X15Y135_SLICE_X20Y135_BO6;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C = CLBLM_R_X15Y135_SLICE_X20Y135_CO6;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D = CLBLM_R_X15Y135_SLICE_X20Y135_DO6;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_AMUX = CLBLM_R_X15Y135_SLICE_X20Y135_A_XOR;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_BMUX = CLBLM_R_X15Y135_SLICE_X20Y135_B_XOR;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_CMUX = CLBLM_R_X15Y135_SLICE_X20Y135_C_XOR;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_DMUX = CLBLM_R_X15Y135_SLICE_X20Y135_D_XOR;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A = CLBLM_R_X15Y135_SLICE_X21Y135_AO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B = CLBLM_R_X15Y135_SLICE_X21Y135_BO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C = CLBLM_R_X15Y135_SLICE_X21Y135_CO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D = CLBLM_R_X15Y135_SLICE_X21Y135_DO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_DMUX = CLBLM_R_X15Y135_SLICE_X21Y135_DO5;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_A = CLBLM_R_X15Y136_SLICE_X20Y136_AO6;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_B = CLBLM_R_X15Y136_SLICE_X20Y136_BO6;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_C = CLBLM_R_X15Y136_SLICE_X20Y136_CO6;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_D = CLBLM_R_X15Y136_SLICE_X20Y136_DO6;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_AMUX = CLBLM_R_X15Y136_SLICE_X20Y136_A_XOR;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_BMUX = CLBLM_R_X15Y136_SLICE_X20Y136_B_XOR;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_CMUX = CLBLM_R_X15Y136_SLICE_X20Y136_C_XOR;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_DMUX = CLBLM_R_X15Y136_SLICE_X20Y136_D_XOR;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_A = CLBLM_R_X15Y136_SLICE_X21Y136_AO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_B = CLBLM_R_X15Y136_SLICE_X21Y136_BO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_C = CLBLM_R_X15Y136_SLICE_X21Y136_CO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_D = CLBLM_R_X15Y136_SLICE_X21Y136_DO6;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_A = CLBLM_R_X15Y137_SLICE_X20Y137_AO6;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_B = CLBLM_R_X15Y137_SLICE_X20Y137_BO6;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_C = CLBLM_R_X15Y137_SLICE_X20Y137_CO6;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_D = CLBLM_R_X15Y137_SLICE_X20Y137_DO6;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_AMUX = CLBLM_R_X15Y137_SLICE_X20Y137_A_XOR;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_BMUX = CLBLM_R_X15Y137_SLICE_X20Y137_B_XOR;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_CMUX = CLBLM_R_X15Y137_SLICE_X20Y137_C_XOR;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_DMUX = CLBLM_R_X15Y137_SLICE_X20Y137_D_CY;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_A = CLBLM_R_X15Y137_SLICE_X21Y137_AO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_B = CLBLM_R_X15Y137_SLICE_X21Y137_BO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_C = CLBLM_R_X15Y137_SLICE_X21Y137_CO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_D = CLBLM_R_X15Y137_SLICE_X21Y137_DO6;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_A = CLBLM_R_X15Y138_SLICE_X20Y138_AO6;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_B = CLBLM_R_X15Y138_SLICE_X20Y138_BO6;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_C = CLBLM_R_X15Y138_SLICE_X20Y138_CO6;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_D = CLBLM_R_X15Y138_SLICE_X20Y138_DO6;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_A = CLBLM_R_X15Y138_SLICE_X21Y138_AO6;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_B = CLBLM_R_X15Y138_SLICE_X21Y138_BO6;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_C = CLBLM_R_X15Y138_SLICE_X21Y138_CO6;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_D = CLBLM_R_X15Y138_SLICE_X21Y138_DO6;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_A = CLBLM_R_X15Y139_SLICE_X20Y139_AO6;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_B = CLBLM_R_X15Y139_SLICE_X20Y139_BO6;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_C = CLBLM_R_X15Y139_SLICE_X20Y139_CO6;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_D = CLBLM_R_X15Y139_SLICE_X20Y139_DO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_A = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_B = CLBLM_R_X15Y139_SLICE_X21Y139_BO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_C = CLBLM_R_X15Y139_SLICE_X21Y139_CO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_D = CLBLM_R_X15Y139_SLICE_X21Y139_DO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_AMUX = CLBLM_R_X15Y139_SLICE_X21Y139_AO5;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_BMUX = CLBLM_R_X15Y139_SLICE_X21Y139_BO6;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_A = CLBLM_R_X15Y140_SLICE_X20Y140_AO6;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_B = CLBLM_R_X15Y140_SLICE_X20Y140_BO6;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_C = CLBLM_R_X15Y140_SLICE_X20Y140_CO6;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_D = CLBLM_R_X15Y140_SLICE_X20Y140_DO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_A = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_B = CLBLM_R_X15Y140_SLICE_X21Y140_BO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_C = CLBLM_R_X15Y140_SLICE_X21Y140_CO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_D = CLBLM_R_X15Y140_SLICE_X21Y140_DO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_AMUX = CLBLM_R_X15Y140_SLICE_X21Y140_AO5;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_CMUX = CLBLM_R_X15Y140_SLICE_X21Y140_CO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_A = CLBLM_R_X15Y141_SLICE_X20Y141_AO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_B = CLBLM_R_X15Y141_SLICE_X20Y141_BO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_C = CLBLM_R_X15Y141_SLICE_X20Y141_CO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_D = CLBLM_R_X15Y141_SLICE_X20Y141_DO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_A = CLBLM_R_X15Y141_SLICE_X21Y141_AO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_B = CLBLM_R_X15Y141_SLICE_X21Y141_BO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_C = CLBLM_R_X15Y141_SLICE_X21Y141_CO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_D = CLBLM_R_X15Y141_SLICE_X21Y141_DO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_AMUX = CLBLM_R_X15Y141_SLICE_X21Y141_A5Q;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B = CLBLM_R_X15Y142_SLICE_X20Y142_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C = CLBLM_R_X15Y142_SLICE_X20Y142_CO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_AMUX = CLBLM_R_X15Y142_SLICE_X20Y142_AO5;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_BMUX = CLBLM_R_X15Y142_SLICE_X20Y142_BO5;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_CMUX = CLBLM_R_X15Y142_SLICE_X20Y142_C5Q;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A = CLBLM_R_X15Y142_SLICE_X21Y142_AO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B = CLBLM_R_X15Y142_SLICE_X21Y142_BO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C = CLBLM_R_X15Y142_SLICE_X21Y142_CO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D = CLBLM_R_X15Y142_SLICE_X21Y142_DO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_AMUX = CLBLM_R_X15Y142_SLICE_X21Y142_A5Q;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_CMUX = CLBLM_R_X15Y142_SLICE_X21Y142_CO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_DMUX = CLBLM_R_X15Y142_SLICE_X21Y142_DO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_A = CLBLM_R_X15Y143_SLICE_X20Y143_AO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_B = CLBLM_R_X15Y143_SLICE_X20Y143_BO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_C = CLBLM_R_X15Y143_SLICE_X20Y143_CO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_D = CLBLM_R_X15Y143_SLICE_X20Y143_DO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_AMUX = CLBLM_R_X15Y143_SLICE_X20Y143_AO5;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_A = CLBLM_R_X15Y143_SLICE_X21Y143_AO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_B = CLBLM_R_X15Y143_SLICE_X21Y143_BO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_C = CLBLM_R_X15Y143_SLICE_X21Y143_CO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_D = CLBLM_R_X15Y143_SLICE_X21Y143_DO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_AMUX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_BMUX = CLBLM_R_X15Y143_SLICE_X21Y143_B5Q;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_CMUX = CLBLM_R_X15Y143_SLICE_X21Y143_CO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A = CLBLM_R_X15Y144_SLICE_X20Y144_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B = CLBLM_R_X15Y144_SLICE_X20Y144_BO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D = CLBLM_R_X15Y144_SLICE_X20Y144_DO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_AMUX = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C = CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D = CLBLM_R_X15Y144_SLICE_X21Y144_DO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_A = CLBLM_R_X15Y145_SLICE_X20Y145_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_B = CLBLM_R_X15Y145_SLICE_X20Y145_BO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_C = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_D = CLBLM_R_X15Y145_SLICE_X20Y145_DO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_AMUX = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_A = CLBLM_R_X15Y145_SLICE_X21Y145_AO6;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_B = CLBLM_R_X15Y145_SLICE_X21Y145_BO6;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_C = CLBLM_R_X15Y145_SLICE_X21Y145_CO6;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_D = CLBLM_R_X15Y145_SLICE_X21Y145_DO6;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_A = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_B = CLBLM_R_X15Y146_SLICE_X20Y146_BO6;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_C = CLBLM_R_X15Y146_SLICE_X20Y146_CO6;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_D = CLBLM_R_X15Y146_SLICE_X20Y146_DO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_A = CLBLM_R_X15Y146_SLICE_X21Y146_AO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_B = CLBLM_R_X15Y146_SLICE_X21Y146_BO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_C = CLBLM_R_X15Y146_SLICE_X21Y146_CO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_D = CLBLM_R_X15Y146_SLICE_X21Y146_DO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_AMUX = CLBLM_R_X15Y146_SLICE_X21Y146_F7AMUX_O;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_CMUX = CLBLM_R_X15Y146_SLICE_X21Y146_CO6;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_A = CLBLM_R_X15Y147_SLICE_X20Y147_AO6;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_B = CLBLM_R_X15Y147_SLICE_X20Y147_BO6;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_C = CLBLM_R_X15Y147_SLICE_X20Y147_CO6;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_D = CLBLM_R_X15Y147_SLICE_X20Y147_DO6;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_A = CLBLM_R_X15Y147_SLICE_X21Y147_AO6;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_B = CLBLM_R_X15Y147_SLICE_X21Y147_BO6;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_C = CLBLM_R_X15Y147_SLICE_X21Y147_CO6;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_D = CLBLM_R_X15Y147_SLICE_X21Y147_DO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_A = CLBLM_R_X15Y148_SLICE_X20Y148_AO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_B = CLBLM_R_X15Y148_SLICE_X20Y148_BO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_C = CLBLM_R_X15Y148_SLICE_X20Y148_CO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_D = CLBLM_R_X15Y148_SLICE_X20Y148_DO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_BMUX = CLBLM_R_X15Y148_SLICE_X20Y148_BO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_A = CLBLM_R_X15Y148_SLICE_X21Y148_AO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_B = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_C = CLBLM_R_X15Y148_SLICE_X21Y148_CO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_D = CLBLM_R_X15Y148_SLICE_X21Y148_DO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_AMUX = CLBLM_R_X15Y148_SLICE_X21Y148_AO5;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_A = CLBLM_R_X15Y149_SLICE_X20Y149_AO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_B = CLBLM_R_X15Y149_SLICE_X20Y149_BO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_C = CLBLM_R_X15Y149_SLICE_X20Y149_CO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_D = CLBLM_R_X15Y149_SLICE_X20Y149_DO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_AMUX = CLBLM_R_X15Y149_SLICE_X20Y149_AO5;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_BMUX = CLBLM_R_X15Y149_SLICE_X20Y149_BO5;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_A = CLBLM_R_X15Y149_SLICE_X21Y149_AO6;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_B = CLBLM_R_X15Y149_SLICE_X21Y149_BO6;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_C = CLBLM_R_X15Y149_SLICE_X21Y149_CO6;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_D = CLBLM_R_X15Y149_SLICE_X21Y149_DO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_A = CLBLM_R_X15Y150_SLICE_X20Y150_AO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_B = CLBLM_R_X15Y150_SLICE_X20Y150_BO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_C = CLBLM_R_X15Y150_SLICE_X20Y150_CO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_D = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_DMUX = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_A = CLBLM_R_X15Y150_SLICE_X21Y150_AO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_B = CLBLM_R_X15Y150_SLICE_X21Y150_BO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_C = CLBLM_R_X15Y150_SLICE_X21Y150_CO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_D = CLBLM_R_X15Y150_SLICE_X21Y150_DO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_AMUX = CLBLM_R_X15Y150_SLICE_X21Y150_AO5;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_CMUX = CLBLM_R_X15Y150_SLICE_X21Y150_CO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A = CLBLM_R_X15Y151_SLICE_X20Y151_AO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B = CLBLM_R_X15Y151_SLICE_X20Y151_BO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C = CLBLM_R_X15Y151_SLICE_X20Y151_CO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_AMUX = CLBLM_R_X15Y151_SLICE_X20Y151_AO5;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_BMUX = CLBLM_R_X15Y151_SLICE_X20Y151_BO5;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_CMUX = CLBLM_R_X15Y151_SLICE_X20Y151_CO5;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A = CLBLM_R_X15Y151_SLICE_X21Y151_AO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B = CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C = CLBLM_R_X15Y151_SLICE_X21Y151_CO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D = CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_AMUX = CLBLM_R_X15Y151_SLICE_X21Y151_A5Q;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_BMUX = CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_A = CLBLM_R_X15Y152_SLICE_X20Y152_AO6;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_B = CLBLM_R_X15Y152_SLICE_X20Y152_BO6;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_C = CLBLM_R_X15Y152_SLICE_X20Y152_CO6;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_D = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_A = CLBLM_R_X15Y152_SLICE_X21Y152_AO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_B = CLBLM_R_X15Y152_SLICE_X21Y152_BO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_C = CLBLM_R_X15Y152_SLICE_X21Y152_CO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_D = CLBLM_R_X15Y152_SLICE_X21Y152_DO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_AMUX = CLBLM_R_X15Y152_SLICE_X21Y152_AO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_CMUX = CLBLM_R_X15Y152_SLICE_X21Y152_CO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_DMUX = CLBLM_R_X15Y152_SLICE_X21Y152_DO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A = CLBLM_R_X15Y153_SLICE_X20Y153_AO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B = CLBLM_R_X15Y153_SLICE_X20Y153_BO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C = CLBLM_R_X15Y153_SLICE_X20Y153_CO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D = CLBLM_R_X15Y153_SLICE_X20Y153_DO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A = CLBLM_R_X15Y153_SLICE_X21Y153_AO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B = CLBLM_R_X15Y153_SLICE_X21Y153_BO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C = CLBLM_R_X15Y153_SLICE_X21Y153_CO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D = CLBLM_R_X15Y153_SLICE_X21Y153_DO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_AMUX = CLBLM_R_X15Y153_SLICE_X21Y153_AO5;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_CMUX = CLBLM_R_X15Y153_SLICE_X21Y153_CO6;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_OQ = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_TQ = 1'b1;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_OQ = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_TQ = 1'b1;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_OQ = CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_TQ = 1'b1;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_OQ = CLBLL_L_X4Y135_SLICE_X5Y135_B5Q;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_TQ = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_OQ = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_TQ = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_OQ = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_TQ = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_OQ = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_TQ = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_OQ = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_TQ = 1'b1;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_OQ = CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_TQ = 1'b1;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_OQ = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_TQ = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLL_L_X2Y135_SLICE_X1Y135_A5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X2Y137_SLICE_X0Y137_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X2Y137_SLICE_X1Y137_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X2Y137_SLICE_X1Y137_BO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X2Y137_SLICE_X1Y137_AO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y139_SLICE_X1Y139_DO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X2Y137_SLICE_X1Y137_BO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLL_L_X2Y139_SLICE_X1Y139_BO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X2Y139_SLICE_X1Y139_AO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X2Y139_SLICE_X1Y139_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X2Y139_SLICE_X1Y139_BO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X2Y143_SLICE_X0Y143_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X2Y144_SLICE_X0Y144_A5Q;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X2Y147_SLICE_X0Y147_AQ;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_L_X2Y145_SLICE_X0Y145_A5Q;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_O = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_O = LIOB33_X0Y151_IOB_X0Y151_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_O = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_O = LIOB33_X0Y153_IOB_X0Y153_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_O = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_O = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_O = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_O = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_O = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_O = LIOB33_X0Y165_IOB_X0Y166_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_O = LIOB33_X0Y165_IOB_X0Y165_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_O = LIOB33_X0Y167_IOB_X0Y168_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y167_O = LIOB33_X0Y167_IOB_X0Y167_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_O = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_O = LIOB33_X0Y171_IOB_X0Y171_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_O = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_O = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_O = LIOB33_X0Y175_IOB_X0Y176_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_O = LIOB33_X0Y175_IOB_X0Y175_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_O = LIOB33_X0Y177_IOB_X0Y178_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_O = LIOB33_X0Y177_IOB_X0Y177_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_O = LIOB33_X0Y179_IOB_X0Y180_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_O = LIOB33_X0Y179_IOB_X0Y179_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_O = LIOB33_X0Y183_IOB_X0Y184_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_O = LIOB33_X0Y183_IOB_X0Y183_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_O = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_O = LIOB33_X0Y185_IOB_X0Y185_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_O = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_O = LIOB33_X0Y189_IOB_X0Y189_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_O = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_O = LIOB33_X0Y191_IOB_X0Y191_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_O = LIOB33_X0Y195_IOB_X0Y196_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_O = LIOB33_X0Y195_IOB_X0Y195_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_O = LIOB33_X0Y197_IOB_X0Y197_I;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_OQ = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLL_L_X2Y147_SLICE_X0Y147_A5Q;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_O = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign LIOI3_SING_X0Y199_ILOGIC_X0Y199_O = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_OQ = CLBLM_R_X5Y136_SLICE_X7Y136_DQ;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_OQ = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X4Y135_SLICE_X5Y135_A5Q;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLL_L_X2Y139_SLICE_X1Y139_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X2Y139_SLICE_X1Y139_DO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLL_L_X2Y144_SLICE_X0Y144_BQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X2Y144_SLICE_X0Y144_AQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O = LIOB33_X0Y157_IOB_X0Y157_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O = LIOB33_X0Y169_IOB_X0Y170_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O = LIOB33_X0Y169_IOB_X0Y169_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O = LIOB33_X0Y181_IOB_X0Y182_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O = LIOB33_X0Y181_IOB_X0Y181_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O = LIOB33_X0Y193_IOB_X0Y194_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O = LIOB33_X0Y193_IOB_X0Y193_I;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_OQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLL_L_X4Y135_SLICE_X4Y135_C5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X2Y139_SLICE_X1Y139_CO5;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O = LIOB33_X0Y163_IOB_X0Y164_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O = LIOB33_X0Y163_IOB_X0Y163_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O = LIOB33_X0Y187_IOB_X0Y188_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O = LIOB33_X0Y187_IOB_X0Y187_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_OQ = CLBLM_L_X16Y133_SLICE_X23Y133_AQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_OQ = CLBLM_L_X16Y133_SLICE_X23Y133_BQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_OQ = CLBLM_L_X16Y133_SLICE_X22Y133_AQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_TQ = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = CLBLM_L_X16Y133_SLICE_X22Y133_BQ;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = CLBLM_L_X16Y134_SLICE_X23Y134_AQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = CLBLM_L_X16Y133_SLICE_X23Y133_CQ;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = CLBLM_L_X16Y134_SLICE_X22Y134_BQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = CLBLM_L_X16Y135_SLICE_X23Y135_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = CLBLM_L_X16Y139_SLICE_X22Y139_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = CLBLM_L_X16Y138_SLICE_X23Y138_AQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = CLBLM_R_X13Y138_SLICE_X19Y138_BQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = CLBLM_R_X13Y138_SLICE_X19Y138_AQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_OQ = CLBLM_L_X16Y137_SLICE_X23Y137_BQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = CLBLM_L_X16Y138_SLICE_X22Y138_AQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_OQ = CLBLM_L_X16Y139_SLICE_X22Y139_BQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_OQ = CLBLM_L_X16Y137_SLICE_X23Y137_CQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = CLBLM_L_X16Y133_SLICE_X22Y133_CQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = CLBLM_L_X16Y133_SLICE_X23Y133_DQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = CLBLM_R_X13Y138_SLICE_X19Y138_CQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = CLBLM_L_X16Y136_SLICE_X23Y136_DQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = CLBLM_L_X16Y136_SLICE_X23Y136_CQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = CLBLM_L_X16Y136_SLICE_X23Y136_BQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y139_SLICE_X1Y139_DO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X2Y147_SLICE_X0Y147_AQ;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_L_X2Y145_SLICE_X0Y145_A5Q;
  assign RIOB33_SING_X105Y149_IOB_X1Y149_O = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A1 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A2 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A3 = CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A4 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A4 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A5 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A6 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_AX = CLBLL_L_X4Y151_SLICE_X4Y151_DO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_AX = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B4 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B3 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B4 = CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B6 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C4 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C6 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_CE = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C6 = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_CX = CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D1 = CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D4 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A1 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A2 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A3 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A4 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A5 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A6 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = CLBLM_L_X16Y138_SLICE_X23Y138_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_AX = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B2 = CLBLM_R_X7Y139_SLICE_X9Y139_CQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B3 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B5 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B6 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_BX = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C1 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C2 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C3 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A4 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C6 = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CIN = CLBLM_R_X7Y138_SLICE_X8Y138_COUT;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CX = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B4 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D1 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D2 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D3 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C4 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_DX = 1'b0;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D4 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A1 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A3 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A4 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A5 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A6 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_AX = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B1 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B2 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B3 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B4 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B5 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B6 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C1 = CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C2 = CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C3 = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C5 = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C6 = CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A4 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D1 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D2 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D3 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D4 = CLBLM_R_X7Y140_SLICE_X9Y140_F7AMUX_O;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D5 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D6 = CLBLM_R_X7Y137_SLICE_X8Y137_F7AMUX_O;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A2 = CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A3 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A4 = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A5 = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A6 = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B1 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B5 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B6 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C1 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C2 = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C3 = CLBLM_R_X11Y137_SLICE_X15Y137_AO5;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C4 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C5 = CLBLM_R_X7Y141_SLICE_X8Y141_F7AMUX_O;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C6 = CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D2 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D3 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D5 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D6 = CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A4 = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A5 = CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A6 = CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_AX = CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B2 = CLBLM_R_X7Y139_SLICE_X9Y139_CQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B6 = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C1 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C2 = CLBLM_R_X7Y139_SLICE_X9Y139_CQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C3 = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C4 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C5 = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C6 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D1 = CLBLM_R_X7Y139_SLICE_X9Y139_CQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D2 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D3 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D4 = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D6 = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A1 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A3 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A4 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A5 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A6 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_AX = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B1 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B2 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B3 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B4 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B5 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B6 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C2 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C3 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C6 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D1 = CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D2 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D3 = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D4 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D5 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D6 = CLBLM_R_X15Y142_SLICE_X20Y142_AO5;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = CLBLM_R_X13Y138_SLICE_X19Y138_BQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = CLBLM_R_X13Y138_SLICE_X19Y138_AQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A2 = CLBLM_R_X3Y159_SLICE_X3Y159_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A3 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A4 = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A5 = CLBLM_R_X3Y159_SLICE_X2Y159_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B1 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B2 = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B3 = CLBLL_L_X4Y156_SLICE_X4Y156_AO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B4 = CLBLM_R_X3Y157_SLICE_X3Y157_BQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B5 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B6 = CLBLL_L_X2Y158_SLICE_X1Y158_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A1 = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A2 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A3 = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C1 = CLBLL_L_X4Y156_SLICE_X4Y156_BO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C2 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C5 = CLBLL_L_X2Y158_SLICE_X0Y158_A5Q;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C6 = CLBLM_R_X3Y157_SLICE_X3Y157_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_AX = CLBLM_R_X15Y139_SLICE_X21Y139_AO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B2 = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B3 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B6 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C6 = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D3 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D6 = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A3 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_AX = CLBLM_R_X15Y140_SLICE_X21Y140_AO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B2 = CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A2 = CLBLL_L_X4Y156_SLICE_X4Y156_BQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A3 = CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A4 = CLBLL_L_X4Y156_SLICE_X4Y156_CQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A5 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A6 = CLBLM_R_X3Y156_SLICE_X2Y156_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_AX = CLBLL_L_X2Y158_SLICE_X1Y158_CQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B2 = CLBLL_L_X4Y156_SLICE_X4Y156_BQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B3 = CLBLL_L_X2Y158_SLICE_X1Y158_CQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B4 = CLBLL_L_X4Y156_SLICE_X4Y156_CQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B5 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B6 = CLBLM_R_X3Y156_SLICE_X2Y156_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A2 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_BX = CLBLM_R_X3Y157_SLICE_X3Y157_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C1 = CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C2 = CLBLL_L_X4Y156_SLICE_X4Y156_DO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C3 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C4 = CLBLL_L_X2Y158_SLICE_X1Y158_CQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C5 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C6 = CLBLM_R_X3Y156_SLICE_X2Y156_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A4 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A6 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B1 = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_CX = CLBLL_L_X2Y158_SLICE_X0Y158_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D1 = CLBLL_L_X4Y156_SLICE_X4Y156_BQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D2 = CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D3 = CLBLL_L_X4Y156_SLICE_X4Y156_DQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D4 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D5 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D6 = CLBLL_L_X4Y156_SLICE_X4Y156_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_DX = CLBLM_R_X3Y156_SLICE_X2Y156_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A1 = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A2 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A4 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A5 = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A6 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B4 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B6 = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CE = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D3 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D4 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D5 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_D1 = CLBLM_L_X16Y137_SLICE_X23Y137_BQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_T1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = CLBLM_L_X16Y138_SLICE_X22Y138_AQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y63_T1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A1 = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A2 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A4 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A5 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A6 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_AX = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B1 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B4 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B6 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_BX = CLBLM_R_X15Y143_SLICE_X21Y143_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C1 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C2 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C3 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C4 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C5 = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C6 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_CX = CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D1 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D2 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D3 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D4 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D5 = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D6 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A1 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A2 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A3 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A4 = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A5 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A6 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B1 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B2 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B3 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B4 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B6 = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C1 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C2 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C3 = CLBLL_L_X4Y141_SLICE_X5Y141_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C4 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C5 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C6 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D1 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_AO5;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D3 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D4 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D6 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_AX = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B5 = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign LIOB33_X0Y55_IOB_X0Y56_O = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign LIOB33_X0Y55_IOB_X0Y55_O = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C5 = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C6 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_D = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A2 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A3 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A4 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A5 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_AX = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B1 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B2 = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B3 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B5 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B6 = CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C1 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C3 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C4 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C5 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C6 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D2 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D3 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D6 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A1 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A3 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A4 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B1 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B2 = CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B4 = CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C3 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D1 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A3 = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D3 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_AX = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X2Y139_SLICE_X1Y139_CO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C6 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_CE = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D1 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CIN = CLBLM_R_X5Y142_SLICE_X6Y142_COUT;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D3 = CLBLM_R_X3Y141_SLICE_X3Y141_DQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_DX = CLBLM_R_X3Y141_SLICE_X3Y141_DQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D4 = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A6 = CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_AX = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B3 = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D2 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D3 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_D1 = CLBLM_L_X16Y139_SLICE_X22Y139_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A1 = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A3 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A4 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A5 = CLBLM_L_X8Y149_SLICE_X10Y149_CO5;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A6 = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C3 = CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D6 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_T1 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A1 = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A2 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A3 = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A4 = CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A6 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B1 = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B3 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B5 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B6 = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C1 = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C2 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C3 = CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C4 = CLBLM_R_X7Y148_SLICE_X8Y148_CO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C5 = CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D3 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D4 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D6 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_D1 = CLBLM_L_X16Y137_SLICE_X23Y137_CQ;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_T1 = 1'b1;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_D = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_AX = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B4 = CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B6 = CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C2 = CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D1 = CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D3 = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D6 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A1 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B2 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B4 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D1 = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D2 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D3 = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D4 = CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D5 = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D6 = CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_C5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A5 = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A2 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A5 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A2 = CLBLM_R_X5Y151_SLICE_X7Y151_AO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A3 = CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A4 = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B2 = CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A5 = CLBLM_R_X7Y149_SLICE_X8Y149_BO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A6 = CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C1 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B2 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C4 = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C6 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C5 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A2 = CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A3 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A4 = CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A5 = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A6 = CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B4 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C6 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D1 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D2 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D3 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D4 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D5 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A5 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B5 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C1 = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C2 = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C5 = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C6 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B5 = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B6 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_A6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C3 = CLBLM_R_X15Y139_SLICE_X21Y139_AO5;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C4 = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_B6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C5 = CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C6 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_C6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D2 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D4 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X21Y128_D6 = 1'b1;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A1 = CLBLM_R_X15Y128_SLICE_X20Y128_B5Q;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A2 = CLBLM_R_X15Y128_SLICE_X20Y128_BQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A4 = CLBLM_R_X15Y128_SLICE_X20Y128_CQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A5 = CLBLM_R_X15Y128_SLICE_X20Y128_A5Q;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_A6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A2 = CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A5 = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B1 = CLBLM_R_X15Y128_SLICE_X20Y128_B5Q;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B2 = CLBLM_R_X15Y128_SLICE_X20Y128_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B4 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B5 = CLBLM_R_X15Y128_SLICE_X20Y128_A5Q;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C6 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D4 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D2 = CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D3 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D5 = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D6 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D5 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A2 = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A3 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A4 = CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A5 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A6 = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B1 = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B2 = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B3 = CLBLM_L_X16Y142_SLICE_X22Y142_AO5;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C5 = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C6 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D6 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B5 = CLBLM_L_X16Y151_SLICE_X23Y151_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLL_L_X2Y139_SLICE_X1Y139_BO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_DX = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A1 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A2 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A3 = CLBLM_R_X15Y129_SLICE_X21Y129_CQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A4 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A5 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_A6 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B1 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B2 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B3 = CLBLM_R_X15Y129_SLICE_X21Y129_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B5 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_B6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C1 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C2 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C3 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C4 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C5 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_C6 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_CE = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D2 = CLBLM_R_X15Y129_SLICE_X21Y129_CQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D4 = CLBLM_R_X15Y130_SLICE_X21Y130_DO6;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D5 = CLBLM_R_X15Y129_SLICE_X21Y129_AQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_D6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_R_X15Y129_SLICE_X21Y129_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A1 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A2 = CLBLM_R_X15Y129_SLICE_X20Y129_BQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A3 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A4 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A5 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_A6 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A2 = CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A3 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A5 = CLBLM_R_X7Y151_SLICE_X8Y151_BO5;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B1 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B5 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B6 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C4 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C5 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C6 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_CE = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A1 = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A2 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A4 = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B4 = CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A1 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A2 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A3 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A4 = CLBLM_R_X3Y131_SLICE_X2Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A5 = CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A6 = CLBLL_L_X2Y131_SLICE_X1Y131_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D2 = CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D3 = CLBLM_R_X5Y151_SLICE_X6Y151_CO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_AX = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B1 = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B2 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B3 = CLBLM_R_X3Y131_SLICE_X2Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B4 = CLBLL_L_X2Y131_SLICE_X1Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B5 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B6 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_BX = CLBLL_L_X4Y133_SLICE_X5Y133_F7AMUX_O;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C1 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C2 = CLBLM_R_X3Y131_SLICE_X2Y131_CQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C3 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C4 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C6 = CLBLL_L_X2Y131_SLICE_X1Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CE = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CX = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1 = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A1 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A2 = CLBLM_R_X15Y130_SLICE_X21Y130_BQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A3 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A5 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_A6 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B1 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B2 = CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B3 = CLBLM_R_X15Y130_SLICE_X21Y130_CQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B5 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_B6 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C1 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C2 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C3 = CLBLM_L_X16Y131_SLICE_X22Y131_AQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C5 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_C6 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_CE = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D2 = CLBLM_R_X15Y130_SLICE_X21Y130_CQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D3 = CLBLM_L_X16Y131_SLICE_X22Y131_AQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D4 = CLBLM_R_X15Y130_SLICE_X21Y130_BQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D5 = CLBLM_R_X15Y130_SLICE_X21Y130_AQ;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_D6 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X21Y130_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A1 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A2 = CLBLM_R_X13Y136_SLICE_X19Y136_BQ;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A3 = CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A5 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_A6 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_AX = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B2 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_B6 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C2 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_C6 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_CE = CLBLM_R_X15Y130_SLICE_X20Y130_AO6;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D1 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D2 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D3 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D4 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D5 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A6 = 1'b1;
  assign CLBLM_R_X15Y130_SLICE_X20Y130_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A1 = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A2 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A4 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A5 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A6 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B1 = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B2 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B4 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B5 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B6 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C1 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C2 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C3 = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C4 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C5 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C6 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D1 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D2 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D3 = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D4 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D5 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D6 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A1 = CLBLM_R_X15Y129_SLICE_X21Y129_B5Q;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A2 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A3 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A4 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A5 = CLBLM_R_X13Y136_SLICE_X19Y136_AQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_A6 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_AX = CLBLM_R_X15Y131_SLICE_X21Y131_BO5;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B1 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B2 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B3 = CLBLM_R_X15Y131_SLICE_X21Y131_AQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B4 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B5 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_B6 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C1 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C2 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C3 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C4 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C5 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_C6 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_CE = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D1 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D2 = CLBLM_R_X15Y131_SLICE_X21Y131_CQ;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D3 = CLBLM_R_X15Y131_SLICE_X21Y131_A5Q;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D4 = CLBLM_R_X15Y129_SLICE_X21Y129_B5Q;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D5 = CLBLM_R_X15Y131_SLICE_X21Y131_AQ;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_B3 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_D6 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X21Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_B4 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A1 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A2 = CLBLM_R_X15Y131_SLICE_X20Y131_BQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A3 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A4 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A5 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_A6 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B1 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B3 = CLBLM_R_X15Y131_SLICE_X20Y131_CQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B4 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B5 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_B6 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C1 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C3 = CLBLM_R_X15Y131_SLICE_X20Y131_DQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C4 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C5 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_C6 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_CE = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_C1 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_C2 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D1 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D3 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D4 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_C3 = 1'b1;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D5 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_D6 = CLBLM_R_X13Y131_SLICE_X19Y131_BQ;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_C4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A1 = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A2 = CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A3 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A4 = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A5 = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A6 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_AX = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLM_R_X15Y131_SLICE_X20Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B1 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B2 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B3 = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B4 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B5 = CLBLM_R_X3Y133_SLICE_X3Y133_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B6 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C1 = CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C2 = CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C3 = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C4 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C5 = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C6 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D1 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D3 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D4 = CLBLM_R_X3Y133_SLICE_X3Y133_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D5 = CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D6 = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A1 = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A2 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A3 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A4 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A5 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B1 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B2 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B3 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B4 = CLBLL_L_X2Y133_SLICE_X1Y133_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B5 = CLBLL_L_X2Y132_SLICE_X1Y132_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C1 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C2 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C6 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_D6 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A1 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A2 = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A3 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A4 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A5 = CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_A6 = CLBLM_R_X15Y129_SLICE_X21Y129_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B2 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B3 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_B6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C2 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C3 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_C6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D2 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D3 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_D6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X17Y128_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A1 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A2 = CLBLM_R_X15Y129_SLICE_X21Y129_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A3 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A4 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A5 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_A6 = CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B2 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B3 = CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B4 = CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B5 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_B6 = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C2 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C3 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_C6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_CE = CLBLM_L_X12Y128_SLICE_X16Y128_BO6;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D1 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D2 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D3 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D4 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D5 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_D6 = 1'b1;
  assign CLBLM_L_X12Y128_SLICE_X16Y128_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B5 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B6 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A1 = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A2 = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A3 = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A4 = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A5 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B1 = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B2 = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B3 = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B4 = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B5 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B6 = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C1 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C2 = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C3 = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C4 = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C5 = CLBLM_R_X3Y133_SLICE_X2Y133_BO5;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C6 = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_CE = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D1 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D2 = CLBLM_R_X3Y133_SLICE_X2Y133_BO5;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D3 = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D4 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D5 = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D6 = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A1 = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A2 = CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A3 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A4 = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A5 = CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A6 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_AX = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B2 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B3 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C2 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D1 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D2 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D3 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D5 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A1 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A2 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A3 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A4 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A5 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_A6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_AX = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B2 = CLBLM_R_X15Y129_SLICE_X21Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B3 = CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B4 = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B5 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_B6 = CLBLM_L_X12Y129_SLICE_X17Y129_AO5;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C1 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C2 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C3 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C4 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C5 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_C6 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_CE = CLBLM_R_X13Y129_SLICE_X18Y129_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D5 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D1 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D2 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D3 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D4 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D5 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_D6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X17Y129_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A1 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A2 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A3 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A4 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A5 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_A6 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B2 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B3 = CLBLM_R_X13Y128_SLICE_X18Y128_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B4 = CLBLM_L_X12Y129_SLICE_X16Y129_CO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B5 = CLBLM_L_X12Y129_SLICE_X16Y129_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_B6 = CLBLM_L_X12Y129_SLICE_X16Y129_AO5;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C1 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C2 = CLBLM_L_X12Y128_SLICE_X17Y128_AQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C3 = CLBLM_R_X15Y129_SLICE_X21Y129_DO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C4 = CLBLM_R_X15Y129_SLICE_X21Y129_BQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C5 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_C6 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A2 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B1 = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D1 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D2 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D3 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D4 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D5 = 1'b1;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B2 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X12Y129_SLICE_X16Y129_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_A1 = CLBLM_R_X15Y133_SLICE_X21Y133_AQ;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_A2 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_A3 = CLBLM_R_X13Y133_SLICE_X19Y133_AQ;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_A4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_A5 = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_A6 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_B1 = CLBLM_R_X15Y134_SLICE_X20Y134_B_XOR;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_B2 = CLBLM_R_X13Y133_SLICE_X19Y133_BQ;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_B3 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_B4 = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_B5 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_B6 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B5 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C2 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_C1 = CLBLM_R_X15Y134_SLICE_X20Y134_D_XOR;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_C2 = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_C3 = CLBLM_R_X13Y133_SLICE_X19Y133_B5Q;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_C4 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_C5 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_C6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_CE = CLBLM_R_X15Y135_SLICE_X21Y135_DO5;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_D1 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_D2 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_D3 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_D4 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_D5 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_D6 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X21Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_A1 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_A2 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_A3 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_A4 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_A5 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_A6 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_B1 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_B2 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_B3 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_B4 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_B5 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_B6 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_C1 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_C2 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_C3 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_C4 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_C5 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_C6 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_D1 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_D2 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_D3 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_D4 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_D5 = 1'b1;
  assign CLBLM_R_X15Y133_SLICE_X20Y133_D6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A1 = CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A4 = CLBLM_L_X12Y131_SLICE_X17Y131_A5Q;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A5 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_A6 = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_AX = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B1 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B3 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B4 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B5 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_B6 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C2 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C4 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C5 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_C6 = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_CE = CLBLM_R_X13Y130_SLICE_X18Y130_CO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C1 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C2 = CLBLM_R_X15Y153_SLICE_X21Y153_AO6;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D2 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D3 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D4 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D5 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_D6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C3 = CLBLM_L_X16Y150_SLICE_X22Y150_B_XOR;
  assign CLBLM_L_X12Y130_SLICE_X17Y130_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A2 = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A3 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A4 = CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A5 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_A6 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B1 = CLBLM_L_X12Y130_SLICE_X16Y130_DO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B2 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B3 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B4 = CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B5 = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_B6 = CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C1 = CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C2 = CLBLM_L_X12Y130_SLICE_X17Y130_AO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C3 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C4 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C5 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_C6 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_CE = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D3 = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D4 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D5 = CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_D6 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X12Y130_SLICE_X16Y130_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_A1 = CLBLM_R_X15Y134_SLICE_X20Y134_A_XOR;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_A2 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_A3 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_A4 = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_A5 = CLBLM_R_X13Y134_SLICE_X19Y134_AQ;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_A6 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_B1 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_B2 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_B3 = CLBLM_R_X15Y134_SLICE_X20Y134_C_XOR;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_B4 = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_B5 = CLBLM_R_X13Y133_SLICE_X19Y133_A5Q;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_B6 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_C1 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_C2 = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_C3 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_C4 = CLBLM_R_X15Y135_SLICE_X20Y135_A_XOR;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_C5 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_C6 = CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_CE = CLBLM_R_X15Y135_SLICE_X21Y135_DO5;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_D1 = CLBLM_R_X15Y135_SLICE_X21Y135_AQ;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_D2 = CLBLM_R_X15Y136_SLICE_X21Y136_CQ;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_D3 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_D4 = CLBLM_R_X15Y134_SLICE_X21Y134_BQ;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_D5 = CLBLM_R_X15Y134_SLICE_X21Y134_AQ;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_D6 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X21Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_A1 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_A2 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_A3 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_A4 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_A5 = CLBLM_R_X15Y134_SLICE_X21Y134_AQ;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_A6 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_AX = CLBLM_R_X15Y133_SLICE_X21Y133_AQ;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_B1 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_B2 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_B3 = CLBLM_R_X15Y131_SLICE_X20Y131_BQ;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_B4 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_B5 = CLBLM_R_X15Y133_SLICE_X21Y133_BQ;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_B6 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_BX = 1'b0;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_C1 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_C2 = CLBLM_R_X15Y134_SLICE_X21Y134_BQ;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_C3 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_C4 = CLBLM_R_X15Y131_SLICE_X20Y131_CQ;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_C5 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_C6 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_CE = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_CX = 1'b0;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_D1 = CLBLM_R_X15Y133_SLICE_X21Y133_CQ;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_D2 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_D3 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_D4 = CLBLM_R_X15Y131_SLICE_X20Y131_DQ;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_D5 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_D6 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_DX = 1'b0;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A1 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A2 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A6 = 1'b1;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B1 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B2 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C1 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C2 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D1 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D2 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A1 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A2 = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A3 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_AX = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign LIOB33_SING_X0Y50_IOB_X0Y50_O = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B1 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B2 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D = LIOB33_X0Y187_IOB_X0Y188_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_BX = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C1 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C2 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D1 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D2 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A1 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A2 = CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A3 = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A4 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A5 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B1 = CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B2 = CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B3 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B5 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B6 = CLBLM_R_X13Y132_SLICE_X18Y132_AO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C2 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C4 = CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C5 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C6 = CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_CE = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D1 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D5 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D6 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A1 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A2 = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A3 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A4 = CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A5 = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B2 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B4 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B5 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C2 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C4 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C5 = CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C6 = CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_CE = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D3 = CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D4 = CLBLM_L_X12Y130_SLICE_X17Y130_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D5 = CLBLM_L_X12Y132_SLICE_X17Y132_A5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D6 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A1 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A2 = CLBLM_R_X13Y134_SLICE_X19Y134_B5Q;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A3 = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A5 = CLBLM_R_X15Y135_SLICE_X20Y135_B_XOR;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_A6 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B1 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B2 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B3 = CLBLM_R_X15Y135_SLICE_X20Y135_C_XOR;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B4 = CLBLM_R_X13Y134_SLICE_X19Y134_A5Q;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B5 = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_B6 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C1 = CLBLM_R_X15Y136_SLICE_X21Y136_AQ;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C2 = CLBLM_R_X15Y134_SLICE_X21Y134_DO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C3 = CLBLM_R_X15Y138_SLICE_X21Y138_BQ;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C5 = CLBLM_R_X15Y136_SLICE_X21Y136_DQ;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_C6 = CLBLM_R_X15Y137_SLICE_X21Y137_BQ;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_CE = CLBLM_R_X15Y135_SLICE_X21Y135_DO5;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D1 = CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D2 = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D4 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_D6 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X21Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_A6 = CLBLM_R_X15Y134_SLICE_X21Y134_CQ;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_AX = 1'b0;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_B6 = CLBLM_R_X15Y135_SLICE_X21Y135_AQ;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_BX = 1'b0;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_C6 = CLBLM_R_X15Y135_SLICE_X21Y135_BQ;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_CIN = CLBLM_R_X15Y134_SLICE_X20Y134_COUT;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_CX = 1'b0;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D1 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D2 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D3 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D4 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D5 = 1'b1;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_D6 = CLBLM_R_X15Y136_SLICE_X21Y136_AQ;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_DX = 1'b0;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_AX = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_BX = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_CE = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_CX = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_DX = CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A1 = CLBLM_R_X3Y134_SLICE_X3Y134_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A3 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A5 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A6 = CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_AX = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_BX = CLBLM_R_X3Y134_SLICE_X3Y134_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_CE = CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_CX = CLBLM_R_X3Y134_SLICE_X3Y134_CQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A1 = CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A2 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A3 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A4 = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A5 = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_DX = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B1 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B2 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B3 = CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B4 = CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C2 = CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C4 = CLBLM_L_X12Y132_SLICE_X17Y132_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C5 = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C6 = CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_CE = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D1 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D2 = CLBLM_L_X12Y131_SLICE_X17Y131_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D3 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D4 = CLBLM_L_X12Y132_SLICE_X17Y132_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D5 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D6 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A1 = CLBLM_L_X12Y131_SLICE_X17Y131_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A2 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A3 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A4 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A5 = CLBLM_L_X12Y132_SLICE_X17Y132_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B1 = CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B2 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B3 = CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B6 = CLBLM_L_X12Y131_SLICE_X17Y131_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C2 = CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C4 = CLBLM_L_X12Y132_SLICE_X16Y132_AO5;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C5 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C6 = CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D3 = CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D4 = CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D5 = CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D6 = CLBLM_L_X12Y132_SLICE_X17Y132_B5Q;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_A1 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_A2 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_A3 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_A4 = CLBLM_R_X15Y135_SLICE_X20Y135_D_XOR;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_A5 = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_A6 = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_B1 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_B2 = CLBLM_R_X13Y136_SLICE_X18Y136_BQ;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_B3 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_B4 = CLBLM_R_X15Y136_SLICE_X20Y136_B_XOR;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_B5 = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_B6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_C1 = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_C2 = CLBLM_R_X13Y136_SLICE_X18Y136_A5Q;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_C3 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_C4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_C5 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_C6 = CLBLM_R_X15Y136_SLICE_X20Y136_C_XOR;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_CE = CLBLM_R_X15Y135_SLICE_X21Y135_DO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_D1 = CLBLM_R_X13Y136_SLICE_X18Y136_B5Q;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_D2 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_D3 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_D4 = CLBLM_R_X15Y136_SLICE_X20Y136_D_XOR;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_D5 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_D6 = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X15Y136_SLICE_X21Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_A1 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_A2 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_A3 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_A4 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_A5 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_A6 = CLBLM_R_X15Y137_SLICE_X21Y137_AQ;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_AX = 1'b0;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLL_L_X2Y135_SLICE_X1Y135_A5Q;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_B1 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_B2 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_B3 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_B4 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_B5 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_B6 = CLBLM_R_X15Y136_SLICE_X21Y136_BQ;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_BX = 1'b0;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_C1 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_C2 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_C3 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_C4 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_C5 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_C6 = CLBLM_R_X15Y136_SLICE_X21Y136_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_CIN = CLBLM_R_X15Y135_SLICE_X20Y135_COUT;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_CX = 1'b0;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_D1 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_D2 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_D3 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_D4 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_D5 = 1'b1;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_D6 = CLBLM_R_X15Y136_SLICE_X21Y136_DQ;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_DX = 1'b0;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A2 = CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A3 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A6 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A1 = CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A3 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A4 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A6 = CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_AX = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B2 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B3 = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B4 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B5 = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B6 = CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C1 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C2 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C5 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C6 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_CE = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D1 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D2 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D5 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D6 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A1 = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A2 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A3 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A4 = CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A5 = CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A6 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B2 = CLBLM_L_X12Y133_SLICE_X16Y133_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B3 = CLBLM_R_X13Y135_SLICE_X19Y135_DQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B4 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B5 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C2 = CLBLM_R_X13Y133_SLICE_X18Y133_BO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C3 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C4 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C5 = CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C6 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D1 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D2 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D3 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D5 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D6 = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_A1 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_A2 = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_A3 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_A4 = CLBLM_R_X13Y138_SLICE_X18Y138_AQ;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_A5 = CLBLM_R_X15Y136_SLICE_X20Y136_A_XOR;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_A6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_B1 = CLBLM_L_X12Y138_SLICE_X17Y138_AQ;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_B2 = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_B3 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_B4 = CLBLM_R_X15Y137_SLICE_X20Y137_A_XOR;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_B5 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_B6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_C1 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_C2 = CLBLL_L_X26Y135_SLICE_X38Y135_AO5;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_C3 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_C5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_C6 = CLBLL_L_X26Y135_SLICE_X38Y135_AO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_CE = CLBLM_R_X15Y135_SLICE_X21Y135_DO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_D1 = CLBLM_R_X15Y134_SLICE_X20Y134_CQ;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_D2 = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_D4 = CLBLM_L_X16Y136_SLICE_X23Y136_AQ;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_D5 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_D6 = CLBLL_L_X26Y135_SLICE_X38Y135_AO6;
  assign CLBLM_R_X15Y137_SLICE_X21Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_A1 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_A2 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_A3 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_A4 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_A5 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_A6 = CLBLM_R_X15Y137_SLICE_X21Y137_BQ;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_AX = 1'b0;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_B1 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_B2 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_B3 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_B4 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_B5 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_B6 = CLBLM_R_X15Y138_SLICE_X21Y138_AQ;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_BX = 1'b0;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_C1 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_C2 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_C3 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_C4 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_C5 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_C6 = CLBLM_R_X15Y138_SLICE_X21Y138_BQ;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_CIN = CLBLM_R_X15Y136_SLICE_X20Y136_COUT;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_CX = 1'b0;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_D1 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_D2 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_D3 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_D4 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_D5 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_D6 = 1'b1;
  assign CLBLM_R_X15Y137_SLICE_X20Y137_DX = 1'b0;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_AX = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_CE = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A1 = CLBLM_R_X3Y126_SLICE_X2Y126_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A2 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A3 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A4 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A5 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B1 = CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B2 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B3 = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B4 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B6 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C1 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C2 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C3 = CLBLM_R_X3Y126_SLICE_X2Y126_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C4 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C5 = CLBLM_R_X15Y137_SLICE_X20Y137_D_CY;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C6 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D1 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D2 = CLBLM_R_X13Y133_SLICE_X18Y133_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D3 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D4 = CLBLM_R_X13Y135_SLICE_X19Y135_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D6 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A1 = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A2 = CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A3 = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A4 = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A6 = CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B1 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B2 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B3 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B4 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B5 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B6 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C2 = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C3 = CLBLM_R_X3Y126_SLICE_X2Y126_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C4 = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C5 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C6 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A2 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D2 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D3 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D4 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D6 = CLBLM_R_X3Y126_SLICE_X2Y126_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A5 = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A6 = CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_A1 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_A2 = CLBLM_R_X15Y137_SLICE_X20Y137_B_XOR;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_A3 = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_A4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_A5 = CLBLM_L_X12Y138_SLICE_X17Y138_BQ;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_A6 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B1 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_B1 = CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_B2 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_B3 = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_B4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_B5 = CLBLM_R_X15Y137_SLICE_X20Y137_C_XOR;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_B6 = CLBLM_R_X13Y138_SLICE_X18Y138_A5Q;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_C1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B4 = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_C2 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_C3 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_C4 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_C5 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_C6 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_CE = CLBLM_R_X15Y135_SLICE_X21Y135_DO6;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_D1 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_D2 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_D3 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_D4 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_D5 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_D6 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X21Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_A1 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_A2 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_A3 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_A4 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_A5 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_A6 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_B1 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_B2 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_B3 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_B4 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_B5 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_B6 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_C1 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_C2 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_C3 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_C4 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_C5 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_C6 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_D1 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_D2 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_D3 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_D4 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_D5 = 1'b1;
  assign CLBLM_R_X15Y138_SLICE_X20Y138_D6 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A1 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A3 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A4 = CLBLM_R_X3Y140_SLICE_X2Y140_BO5;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A6 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_AX = 1'b0;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B1 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B2 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B3 = CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B4 = CLBLL_L_X2Y140_SLICE_X1Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B5 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B6 = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A6 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_BX = CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C1 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C2 = CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C3 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C4 = CLBLL_L_X2Y140_SLICE_X1Y140_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C5 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C6 = CLBLL_L_X2Y140_SLICE_X1Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_CE = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_CX = CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D1 = CLBLL_L_X2Y140_SLICE_X1Y140_CQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D2 = CLBLL_L_X2Y140_SLICE_X1Y140_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D3 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D4 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D5 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D6 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A2 = CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A3 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A4 = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B3 = CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B1 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B2 = CLBLL_L_X2Y140_SLICE_X1Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B3 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B4 = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B5 = CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B5 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B6 = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C1 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C3 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C4 = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D3 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D4 = CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A2 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A3 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A4 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A5 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A6 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_AX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B1 = CLBLM_L_X16Y134_SLICE_X22Y134_AO5;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B3 = CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B4 = CLBLM_L_X12Y137_SLICE_X16Y137_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B5 = CLBLM_R_X15Y134_SLICE_X20Y134_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C1 = CLBLM_R_X3Y126_SLICE_X2Y126_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C2 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C3 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C5 = CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C6 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_CE = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C5 = CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D2 = CLBLM_R_X13Y135_SLICE_X19Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D3 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D4 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D5 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D6 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A1 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A2 = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A3 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A4 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A5 = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B1 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B2 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B4 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B5 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B6 = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C1 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C4 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C6 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D1 = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D3 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D4 = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D6 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D3 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D4 = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D6 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_A1 = CLBLM_R_X15Y139_SLICE_X21Y139_BO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_A2 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_A3 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_A4 = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_A5 = CLBLM_R_X15Y141_SLICE_X21Y141_DO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_A6 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_AX = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_B1 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_B2 = CLBLM_L_X16Y140_SLICE_X22Y140_CQ;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_B3 = CLBLM_R_X15Y140_SLICE_X21Y140_DQ;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_B4 = CLBLM_R_X15Y139_SLICE_X21Y139_CQ;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_B6 = CLBLM_R_X15Y140_SLICE_X20Y140_CQ;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_BX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_C1 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_C2 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_C3 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_C4 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_C5 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_C6 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_CE = CLBLM_R_X15Y141_SLICE_X20Y141_BO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_CX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_D1 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_D2 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_D3 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_D4 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_D5 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_D6 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X21Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_A1 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_A2 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_A3 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_A4 = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_A5 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_A6 = CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_B1 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_B2 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_B3 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_B4 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_B5 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_B6 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_C1 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_C2 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_C3 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_C4 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_C5 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_C6 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_D1 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_D2 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_D3 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_D4 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_D5 = 1'b1;
  assign CLBLM_R_X15Y139_SLICE_X20Y139_D6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A1 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A3 = CLBLL_L_X2Y140_SLICE_X1Y140_CQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A5 = CLBLL_L_X2Y140_SLICE_X1Y140_DQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B5 = CLBLL_L_X2Y140_SLICE_X1Y140_DQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B6 = CLBLL_L_X2Y141_SLICE_X1Y141_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_BX = CLBLL_L_X2Y140_SLICE_X1Y140_DQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C2 = CLBLL_L_X2Y141_SLICE_X1Y141_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C4 = CLBLL_L_X2Y141_SLICE_X1Y141_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_CE = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_CIN = CLBLM_R_X3Y140_SLICE_X3Y140_COUT;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_CX = CLBLL_L_X2Y141_SLICE_X1Y141_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D1 = CLBLL_L_X2Y141_SLICE_X1Y141_CQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D2 = CLBLL_L_X2Y141_SLICE_X1Y141_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_DX = CLBLL_L_X2Y141_SLICE_X1Y141_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A1 = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A4 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B1 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B2 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B3 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B4 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B5 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B6 = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C2 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C4 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C5 = CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C6 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_CE = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D1 = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D4 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D5 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D6 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A1 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A2 = CLBLM_L_X12Y137_SLICE_X17Y137_CO5;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A3 = CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A5 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A6 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B1 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B2 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B3 = CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B4 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B5 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B6 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C1 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C3 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C4 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C5 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D3 = CLBLL_L_X26Y138_SLICE_X38Y138_AO5;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D4 = CLBLM_R_X13Y131_SLICE_X18Y131_DQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D5 = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D6 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A2 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A3 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A4 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A5 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_AX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B1 = CLBLM_R_X15Y137_SLICE_X21Y137_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B2 = CLBLM_L_X12Y136_SLICE_X16Y136_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B3 = CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B4 = CLBLM_R_X15Y134_SLICE_X21Y134_CQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_BX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C2 = CLBLM_L_X12Y136_SLICE_X16Y136_CQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C3 = CLBLM_L_X10Y133_SLICE_X13Y133_AO5;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C5 = CLBLM_R_X15Y138_SLICE_X21Y138_AQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C6 = CLBLM_R_X15Y135_SLICE_X21Y135_AQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_CE = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_CX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D2 = CLBLM_R_X13Y137_SLICE_X18Y137_CO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D3 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D4 = CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D5 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D6 = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C1 = CLBLM_L_X12Y129_SLICE_X17Y129_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X2Y139_SLICE_X1Y139_CO5;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C2 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_A1 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_A2 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_A3 = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_A4 = CLBLM_R_X15Y141_SLICE_X21Y141_CO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_A5 = CLBLM_R_X15Y140_SLICE_X21Y140_CO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_A6 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_AX = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_B1 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_B2 = CLBLM_R_X15Y139_SLICE_X21Y139_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C3 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_B3 = CLBLM_R_X15Y140_SLICE_X21Y140_AQ;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_B4 = CLBLM_L_X16Y140_SLICE_X22Y140_AQ;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_B5 = CLBLM_R_X15Y140_SLICE_X20Y140_AQ;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_BX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_C1 = CLBLM_L_X16Y140_SLICE_X22Y140_BQ;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_C2 = CLBLM_R_X15Y140_SLICE_X21Y140_CQ;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_C3 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_C5 = CLBLM_R_X15Y139_SLICE_X21Y139_BQ;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_C6 = CLBLM_R_X15Y140_SLICE_X20Y140_BQ;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_CE = CLBLM_R_X13Y141_SLICE_X19Y141_AO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_CX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_D1 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_D2 = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C4 = CLBLM_R_X13Y128_SLICE_X18Y128_A5Q;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_D3 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_D4 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_D5 = CLBLM_R_X15Y141_SLICE_X21Y141_BO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_D6 = CLBLM_R_X15Y140_SLICE_X21Y140_BO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_DX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_R_X15Y140_SLICE_X21Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_A1 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_A2 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_A3 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_A4 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_A5 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_A6 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_AX = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_B1 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_B2 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_B3 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_B4 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_B5 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_B6 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_BX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_C1 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_C2 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_C3 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_C4 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_C5 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_C6 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_CE = CLBLM_R_X15Y141_SLICE_X20Y141_AO6;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_CX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_D1 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_D2 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_D3 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_D4 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_D5 = 1'b1;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_D6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A3 = CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A6 = CLBLL_L_X2Y141_SLICE_X1Y141_CQ;
  assign CLBLM_R_X15Y140_SLICE_X20Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_AX = CLBLL_L_X2Y141_SLICE_X1Y141_CQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B2 = CLBLL_L_X2Y142_SLICE_X1Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B3 = CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_BX = CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C2 = CLBLL_L_X2Y142_SLICE_X1Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C4 = CLBLL_L_X2Y142_SLICE_X1Y142_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_CE = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_CIN = CLBLM_R_X3Y141_SLICE_X3Y141_COUT;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_CX = CLBLL_L_X2Y142_SLICE_X1Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D3 = CLBLL_L_X2Y142_SLICE_X1Y142_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D5 = CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_DX = CLBLL_L_X2Y142_SLICE_X1Y142_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A1 = CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A2 = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A4 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_AX = CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B2 = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B4 = CLBLL_L_X4Y141_SLICE_X5Y141_CQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B5 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B6 = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C1 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C2 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C3 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C4 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C6 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D1 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D2 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D3 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D4 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D5 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D6 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign RIOB33_X105Y125_IOB_X1Y126_O = CLBLM_L_X16Y133_SLICE_X23Y133_BQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A2 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A3 = CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A4 = CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A6 = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B2 = CLBLM_L_X12Y137_SLICE_X17Y137_BQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B3 = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B4 = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B5 = CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B6 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C1 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C2 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C3 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C4 = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C5 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D1 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D2 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D3 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D4 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D5 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D6 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A1 = CLBLM_R_X13Y138_SLICE_X19Y138_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A3 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B2 = CLBLM_L_X12Y137_SLICE_X16Y137_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B3 = CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B4 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B5 = CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B6 = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C1 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C2 = CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C4 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C5 = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X2Y137_SLICE_X0Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D1 = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D3 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D6 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_A1 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_A2 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_A3 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_A4 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_A5 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_A6 = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_AX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_B1 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_B3 = CLBLM_R_X15Y141_SLICE_X21Y141_AQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_B4 = CLBLM_R_X15Y141_SLICE_X20Y141_BQ;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_A4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_B5 = CLBLM_L_X16Y141_SLICE_X23Y141_AQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_B6 = CLBLM_R_X15Y142_SLICE_X21Y142_CQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_BX = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_C1 = CLBLM_L_X16Y141_SLICE_X22Y141_BQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_C2 = CLBLM_R_X15Y141_SLICE_X20Y141_DQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_C3 = CLBLM_R_X15Y141_SLICE_X21Y141_DQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_C4 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_C5 = CLBLM_L_X16Y141_SLICE_X23Y141_CQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_CE = CLBLM_R_X15Y141_SLICE_X20Y141_CO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_CX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_D1 = CLBLM_L_X16Y141_SLICE_X23Y141_DQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_D2 = CLBLM_R_X13Y141_SLICE_X19Y141_CQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_D3 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_D4 = CLBLM_R_X15Y141_SLICE_X21Y141_A5Q;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_D5 = CLBLM_L_X16Y141_SLICE_X22Y141_CQ;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_DX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_R_X15Y141_SLICE_X21Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_A1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_A2 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_B1 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_A3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_A4 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_B2 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_AX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_B1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_B2 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_B5 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_B4 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_BX = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_C1 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_C2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_C3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_C5 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_C6 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_CE = CLBLM_L_X16Y141_SLICE_X22Y141_AO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_D1 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_CX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_D1 = CLBLM_R_X15Y143_SLICE_X21Y143_DO6;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_D2 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_D2 = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_D4 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_D5 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_D6 = CLBLM_L_X16Y141_SLICE_X22Y141_CO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_D3 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_DX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A3 = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A5 = CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A6 = 1'b1;
  assign CLBLM_R_X15Y141_SLICE_X20Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_AX = CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B2 = CLBLL_L_X2Y143_SLICE_X1Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B3 = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_BX = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C2 = CLBLL_L_X2Y143_SLICE_X1Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C4 = CLBLL_L_X2Y143_SLICE_X1Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CE = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CIN = CLBLM_R_X3Y142_SLICE_X3Y142_COUT;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_C6 = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CX = CLBLL_L_X2Y143_SLICE_X1Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D1 = CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D2 = CLBLL_L_X2Y143_SLICE_X1Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_DX = 1'b0;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D3 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A2 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A3 = CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A5 = CLBLL_L_X4Y141_SLICE_X5Y141_BQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A6 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B2 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B3 = CLBLL_L_X4Y141_SLICE_X5Y141_DQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B5 = CLBLL_L_X2Y158_SLICE_X0Y158_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B6 = CLBLM_R_X3Y137_SLICE_X2Y137_CQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C1 = CLBLM_R_X3Y137_SLICE_X2Y137_DQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C2 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C3 = CLBLM_R_X3Y158_SLICE_X2Y158_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C4 = CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_D1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D2 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D3 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D4 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D6 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A2 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A3 = CLBLM_L_X12Y137_SLICE_X17Y137_BQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A4 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A5 = CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A6 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_AX = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B1 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B2 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B3 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_BX = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C1 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C2 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C3 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C6 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_CE = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D1 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D2 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D3 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D6 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_BI = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_CE = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_DI = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A1 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A2 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A6 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_AX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B1 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B2 = CLBLM_R_X15Y142_SLICE_X21Y142_BQ;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B3 = CLBLM_R_X15Y141_SLICE_X20Y141_AQ;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B4 = CLBLM_R_X15Y144_SLICE_X21Y144_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B6 = CLBLM_L_X16Y142_SLICE_X22Y142_BQ;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_BX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D6 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C1 = CLBLM_R_X13Y141_SLICE_X19Y141_BQ;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C2 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C3 = CLBLM_R_X15Y144_SLICE_X21Y144_CQ;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C4 = CLBLM_R_X15Y142_SLICE_X21Y142_A5Q;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C6 = CLBLM_L_X16Y142_SLICE_X22Y142_DQ;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_CE = CLBLM_L_X16Y141_SLICE_X22Y141_BO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_CX = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D1 = CLBLM_R_X15Y140_SLICE_X21Y140_BQ;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D2 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D3 = CLBLM_R_X15Y143_SLICE_X21Y143_B5Q;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D4 = CLBLM_L_X16Y143_SLICE_X22Y143_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D5 = CLBLM_R_X15Y142_SLICE_X20Y142_C5Q;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_DX = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C1 = CLBLM_L_X16Y152_SLICE_X22Y152_D_XOR;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A1 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A2 = CLBLM_R_X15Y142_SLICE_X21Y142_DO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A3 = CLBLM_R_X15Y142_SLICE_X21Y142_CO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A4 = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A5 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A6 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_C3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_AX = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_C4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B1 = CLBLM_R_X15Y143_SLICE_X20Y143_CO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B2 = CLBLM_L_X16Y142_SLICE_X22Y142_DO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B3 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B4 = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_C5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B5 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C2 = CLBLM_R_X15Y150_SLICE_X21Y150_CO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_BX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C1 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C2 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C6 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_CE = CLBLM_R_X15Y141_SLICE_X20Y141_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_CX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D1 = CLBLM_L_X16Y142_SLICE_X22Y142_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D2 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D4 = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D5 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D6 = CLBLM_R_X15Y143_SLICE_X20Y143_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_DX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A1 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A2 = CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A3 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A4 = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A5 = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A6 = CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_AX = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B1 = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B2 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B3 = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B4 = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B5 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B6 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C1 = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C2 = CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C3 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C5 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C6 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_D1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_D2 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_D3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D1 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D2 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D4 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D6 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B5 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C5 = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B6 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A2 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A4 = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C4 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_D6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B1 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B3 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B4 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B5 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B6 = CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C1 = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C2 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C3 = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C4 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C5 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C6 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D2 = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D3 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D4 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D5 = CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D6 = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A3 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A4 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A5 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A6 = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B1 = CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B2 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B3 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B4 = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B5 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B6 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C2 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C3 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C5 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C6 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D1 = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D1 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D2 = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_AI = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_BI = CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A5 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_CE = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_CI = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_DI = 1'b0;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B5 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B6 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_A1 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_A2 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_A3 = CLBLM_R_X15Y142_SLICE_X21Y142_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_A4 = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_A5 = CLBLM_R_X15Y143_SLICE_X21Y143_CO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_A6 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_AX = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_B1 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_B2 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_B3 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_B4 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_B5 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_B6 = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_BX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_C1 = CLBLM_L_X16Y143_SLICE_X22Y143_AQ;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_C3 = CLBLM_R_X15Y143_SLICE_X21Y143_BQ;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_C4 = CLBLM_R_X15Y142_SLICE_X20Y142_BQ;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_C5 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_C6 = CLBLM_R_X15Y143_SLICE_X20Y143_BQ;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_CE = CLBLM_R_X15Y141_SLICE_X20Y141_AO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C1 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_CX = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_D1 = CLBLM_L_X16Y143_SLICE_X22Y143_BQ;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_D2 = CLBLM_R_X15Y142_SLICE_X20Y142_DQ;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_D3 = CLBLM_R_X15Y143_SLICE_X21Y143_DQ;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_D4 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_D5 = CLBLM_R_X15Y143_SLICE_X20Y143_DQ;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_DX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_R_X15Y143_SLICE_X21Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_A1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_A2 = CLBLM_R_X15Y144_SLICE_X20Y144_BQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_A3 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_A5 = CLBLM_R_X15Y143_SLICE_X21Y143_AQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_A6 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_AX = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_B1 = CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_B2 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_B3 = CLBLM_R_X15Y143_SLICE_X20Y143_AQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_B4 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_B5 = CLBLM_R_X15Y143_SLICE_X20Y143_AO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X2Y137_SLICE_X1Y137_AO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_BX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_C1 = CLBLM_R_X15Y143_SLICE_X21Y143_AQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_C2 = CLBLM_R_X15Y143_SLICE_X20Y143_AQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_C3 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_C5 = CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_C6 = CLBLM_R_X15Y144_SLICE_X20Y144_BQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_CE = CLBLM_R_X13Y141_SLICE_X19Y141_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_CX = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_D1 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_D2 = CLBLM_R_X15Y143_SLICE_X20Y143_CQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_D3 = CLBLM_R_X15Y142_SLICE_X20Y142_CQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_D4 = CLBLM_R_X15Y143_SLICE_X21Y143_CQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_D5 = CLBLM_R_X15Y144_SLICE_X20Y144_CQ;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_DX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A1 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A2 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A4 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A5 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A6 = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign CLBLM_R_X15Y143_SLICE_X20Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B2 = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B3 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B5 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B6 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A4 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C2 = CLBLM_R_X3Y158_SLICE_X3Y158_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C4 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C5 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C6 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D1 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D2 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D5 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A1 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A4 = CLBLM_R_X3Y140_SLICE_X2Y140_BO5;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A5 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A6 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_AX = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B1 = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B2 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B3 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B4 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B5 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B6 = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A1 = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A2 = CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A3 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A4 = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A5 = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B3 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B1 = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B2 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B5 = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B6 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C1 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C2 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C4 = CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C5 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D1 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D2 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D4 = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D5 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D6 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C5 = CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C6 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C1 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_AI = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C3 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C4 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_BI = CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C5 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_C6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_CI = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_CE = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_DI = 1'b0;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_CIN = CLBLM_L_X16Y153_SLICE_X22Y153_COUT;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A1 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A3 = CLBLM_R_X13Y144_SLICE_X19Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A5 = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_A6 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_AX = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B1 = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B2 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B3 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B4 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B5 = CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_B6 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_BX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C1 = CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C2 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C3 = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C4 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D6 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_C6 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_CE = CLBLM_R_X15Y141_SLICE_X20Y141_CO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_CX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D5 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_D6 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X21Y144_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_DX = 1'b0;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A5 = CLBLM_R_X13Y144_SLICE_X19Y144_CO5;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_A6 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_AX = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B2 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B4 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_B6 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X2Y139_SLICE_X1Y139_AO5;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_BX = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C1 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C2 = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C3 = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C4 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C5 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_C6 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_CE = CLBLM_L_X16Y143_SLICE_X22Y143_AO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_CX = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D1 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D2 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D3 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D4 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D5 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_D6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A1 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A3 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A5 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A6 = 1'b1;
  assign CLBLM_R_X15Y144_SLICE_X20Y144_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B3 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B4 = CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C1 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C2 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C4 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C6 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D1 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D2 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D3 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D4 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A3 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B3 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B4 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B5 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C1 = CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C2 = CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C3 = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C4 = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C5 = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C6 = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D1 = CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D2 = CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D3 = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D4 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D5 = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D6 = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A1 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A2 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A3 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A4 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A5 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_AX = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B2 = CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B3 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B4 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B5 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B6 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C1 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C2 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C3 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C5 = CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C6 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D2 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D4 = CLBLM_L_X12Y141_SLICE_X17Y141_AO5;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D5 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D6 = CLBLM_R_X11Y141_SLICE_X15Y141_CO5;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_AI = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_BI = CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_CE = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_CI = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_DI = 1'b0;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_A1 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_A2 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_A3 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_A4 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_A5 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_A6 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_B1 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_B2 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_B3 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_B4 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_B5 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_B6 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_C1 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_C2 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_C3 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_C4 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_C5 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_C6 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_D1 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_D2 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_D3 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_D4 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_D5 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X21Y145_D6 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_A1 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_A2 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_A3 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_A4 = CLBLM_R_X13Y145_SLICE_X19Y145_BO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_A5 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_A6 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_AX = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_B1 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_B2 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_B3 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_B4 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_B5 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_B6 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_C1 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_C2 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_C3 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_C4 = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_C5 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_C6 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_D1 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_D2 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_D3 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_D4 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_D5 = 1'b1;
  assign CLBLM_R_X15Y145_SLICE_X20Y145_D6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A1 = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A2 = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A4 = CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B1 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B2 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B3 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B6 = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C3 = CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C4 = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C5 = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C6 = CLBLM_R_X15Y143_SLICE_X20Y143_AO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A2 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A3 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A5 = CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B4 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B5 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C2 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C3 = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C6 = CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X2Y137_SLICE_X1Y137_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D1 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D2 = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D3 = CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D5 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A1 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A2 = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A3 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A4 = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A5 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A6 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_AX = CLBLM_R_X15Y142_SLICE_X20Y142_BO5;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B2 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B5 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X2Y137_SLICE_X1Y137_AO5;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C1 = CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C2 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C4 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C5 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C6 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D3 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D4 = CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D5 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D6 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_AI = CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_BI = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_CE = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_CI = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_T1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_DI = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_A1 = CLBLM_R_X15Y146_SLICE_X21Y146_DO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_A2 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_A3 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_A4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_A5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_AX = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_B1 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_B4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_B5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_B6 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_C2 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_C4 = CLBLM_R_X13Y144_SLICE_X19Y144_CO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_C5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_C6 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_A6 = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_D2 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_D3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_D5 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X15Y146_SLICE_X21Y146_D6 = CLBLM_R_X13Y145_SLICE_X19Y145_BO6;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_A1 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_A4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_A5 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_A6 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_A2 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_B1 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_B2 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_B3 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_B4 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_B5 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_B6 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_B2 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_B3 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_C1 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_C2 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_C3 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_C4 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_C5 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_C6 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_D1 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_D2 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_D3 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_D4 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_D5 = 1'b1;
  assign CLBLM_R_X15Y146_SLICE_X20Y146_D6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A1 = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A2 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A3 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A4 = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A6 = CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B1 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B3 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B4 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_C2 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C1 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C5 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_C4 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_C5 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D1 = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D2 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D3 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D4 = CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D5 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D6 = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A1 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A2 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C1 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C2 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C5 = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A1 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A2 = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A3 = CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A5 = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A6 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A1 = CLBLM_L_X12Y137_SLICE_X16Y137_CO5;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A2 = CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A3 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A4 = CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A5 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A6 = CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B1 = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B4 = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B5 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C2 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C3 = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C4 = CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C5 = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C6 = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D1 = CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D6 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_A1 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_A2 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_A4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_B1 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_B2 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_B3 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_B4 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_B5 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_B6 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_C1 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_C2 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_C3 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_C4 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_C5 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_C6 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_D1 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_D2 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_D3 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_D4 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_D5 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X21Y147_D6 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_A1 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_A2 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_A3 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_A4 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_A5 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_A6 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_B1 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_B2 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_B3 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_B4 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_B5 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_B6 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_C1 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_C2 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_C3 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_C4 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_C5 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_C6 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_D1 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_D2 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_D3 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_D4 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_D5 = 1'b1;
  assign CLBLM_R_X15Y147_SLICE_X20Y147_D6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A3 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A4 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A5 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B2 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B5 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C1 = CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C2 = CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C3 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C4 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C6 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D1 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D2 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D3 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D4 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D6 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B1 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B4 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B5 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C1 = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D1 = CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D3 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D4 = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D5 = CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D6 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A2 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A5 = CLBLM_L_X12Y144_SLICE_X17Y144_CO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A6 = CLBLM_R_X13Y145_SLICE_X19Y145_AO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_AX = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B2 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B4 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B5 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C2 = CLBLM_R_X13Y144_SLICE_X18Y144_D_XOR;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C3 = CLBLM_R_X13Y144_SLICE_X18Y144_C_XOR;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C4 = CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C5 = CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D1 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D2 = CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D3 = CLBLM_R_X13Y145_SLICE_X19Y145_BO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D6 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A1 = CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A2 = CLBLM_R_X13Y144_SLICE_X18Y144_B_XOR;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B2 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B5 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C2 = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C3 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C4 = CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C5 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C6 = CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_A6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D5 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_C6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_D6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A3 = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A4 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X2Y137_SLICE_X1Y137_BO5;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_A2 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_A5 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_A6 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_A6 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_B1 = CLBLM_R_X15Y147_SLICE_X21Y147_AO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_B2 = CLBLM_R_X15Y149_SLICE_X21Y149_AO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_B3 = CLBLM_R_X15Y146_SLICE_X21Y146_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_B6 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_C2 = CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_C6 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_D2 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_D3 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C1 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_D4 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_D5 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D1 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D2 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D3 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D4 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D5 = 1'b1;
  assign CLBLL_L_X2Y116_SLICE_X1Y116_D6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C2 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_A1 = CLBLM_R_X15Y148_SLICE_X20Y148_BO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_A2 = CLBLM_R_X15Y150_SLICE_X21Y150_CO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_A3 = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_A4 = CLBLM_L_X16Y152_SLICE_X22Y152_D_XOR;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_A5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_A6 = CLBLM_R_X15Y148_SLICE_X20Y148_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C5 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_B3 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_B4 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_B5 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_B6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_C1 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_C2 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_C3 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_C5 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_C6 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A2 = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_D1 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_D2 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_D3 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_D4 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_D5 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X20Y148_D6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D4 = CLBLM_L_X8Y140_SLICE_X11Y140_AO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A1 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_DQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A3 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_AX = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B1 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B2 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B4 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_BX = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A3 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C2 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C3 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C4 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C5 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C6 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_CE = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A4 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_CX = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D1 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D3 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D4 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D6 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_DX = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A1 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A2 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A3 = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A4 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A5 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B1 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B2 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B3 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B4 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B5 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A5 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C1 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C2 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C3 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C4 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C5 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C6 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A6 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D2 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D3 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D4 = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D5 = CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A1 = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A2 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A4 = CLBLM_R_X13Y148_SLICE_X19Y148_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A5 = CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A6 = CLBLM_R_X15Y149_SLICE_X20Y149_CO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B1 = CLBLM_L_X12Y142_SLICE_X17Y142_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B2 = CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B3 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B4 = CLBLM_R_X13Y148_SLICE_X19Y148_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B5 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B6 = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C1 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C2 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C3 = CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C4 = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C5 = CLBLM_R_X13Y148_SLICE_X19Y148_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C6 = CLBLM_L_X12Y142_SLICE_X17Y142_AO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D2 = CLBLM_R_X13Y145_SLICE_X18Y145_D_XOR;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D4 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D5 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D6 = CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C5 = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A2 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A3 = CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A4 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A5 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B2 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B3 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B4 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B6 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C1 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C2 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C3 = CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C4 = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C5 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C6 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D1 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D2 = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D3 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D4 = CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D5 = CLBLM_R_X13Y148_SLICE_X19Y148_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D6 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X2Y143_SLICE_X0Y143_AQ;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_A1 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_A2 = CLBLM_R_X15Y152_SLICE_X21Y152_BO6;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_A3 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_A5 = CLBLM_R_X15Y149_SLICE_X20Y149_DO6;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_A6 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_B1 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_B2 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_B3 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_B4 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_B5 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_B6 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_C1 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_C2 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_C3 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_C4 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_C5 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_C6 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_D1 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_D2 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_D3 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_D4 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_D5 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X21Y149_D6 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_A1 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_A2 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_A4 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_A6 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_B1 = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_B3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_B4 = CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_B5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_B6 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_C1 = CLBLM_R_X15Y149_SLICE_X20Y149_AO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_C2 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_C3 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_C4 = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_C5 = CLBLM_R_X15Y149_SLICE_X20Y149_BO5;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_C6 = CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_D1 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_D2 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_D3 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_D4 = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_D5 = 1'b1;
  assign CLBLM_R_X15Y149_SLICE_X20Y149_D6 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A1 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A2 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A3 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A4 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A5 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B1 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B3 = CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B4 = CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B5 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B6 = CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C1 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C2 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C3 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C5 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C6 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D1 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D3 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D4 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D5 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A1 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A2 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A3 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A4 = CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A5 = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A6 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B1 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B2 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B3 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B4 = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B5 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B6 = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C1 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C2 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C3 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C4 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C5 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C6 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D1 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D2 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D3 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D4 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D5 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D6 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A2 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A4 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_AX = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B2 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B4 = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B6 = CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C1 = CLBLM_L_X12Y144_SLICE_X17Y144_F7AMUX_O;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C2 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C3 = CLBLM_R_X13Y150_SLICE_X19Y150_F7AMUX_O;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C4 = CLBLM_R_X13Y149_SLICE_X18Y149_F7AMUX_O;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C5 = CLBLM_R_X15Y146_SLICE_X21Y146_F7AMUX_O;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D1 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D2 = CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D4 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D6 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A1 = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A2 = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A3 = CLBLM_R_X15Y148_SLICE_X20Y148_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A4 = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A5 = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A6 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_AX = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B2 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B5 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B6 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C1 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C3 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C4 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C5 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_D = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D1 = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D2 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D3 = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D4 = CLBLM_R_X15Y148_SLICE_X20Y148_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D5 = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D6 = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_A1 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_A2 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_A3 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_A4 = CLBLM_R_X15Y151_SLICE_X21Y151_A5Q;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_A5 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_A6 = 1'b1;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_B2 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_B3 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_B4 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_B5 = CLBLM_L_X16Y152_SLICE_X23Y152_BO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_B6 = CLBLM_R_X15Y149_SLICE_X20Y149_BO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_C1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_C2 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_C4 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_C5 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_C6 = CLBLM_L_X16Y150_SLICE_X22Y150_C_XOR;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_D1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_D2 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_D3 = CLBLM_R_X15Y151_SLICE_X21Y151_A5Q;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_D4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_D5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A6 = 1'b1;
  assign CLBLM_R_X15Y150_SLICE_X21Y150_D6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_AX = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_A1 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B6 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_A2 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_A3 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_BX = 1'b0;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_A4 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C6 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_B1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_B2 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_B3 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_C2 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_CX = 1'b0;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D6 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_C5 = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_C6 = CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_DX = 1'b0;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_D2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A6 = 1'b1;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_D3 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_D4 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A1 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A2 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_AX = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_AX = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B2 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B1 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B2 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B6 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_BX = 1'b0;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C2 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C4 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_CX = 1'b0;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D2 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D4 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D6 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_DX = 1'b0;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A1 = CLBLL_L_X2Y153_SLICE_X0Y153_DQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A2 = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A3 = CLBLM_R_X3Y153_SLICE_X2Y153_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A4 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A5 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A6 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_AX = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B1 = CLBLL_L_X2Y153_SLICE_X0Y153_DQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B2 = CLBLL_L_X2Y153_SLICE_X0Y153_C5Q;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B4 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B6 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C1 = CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C2 = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C3 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C4 = CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_BO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C6 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_CE = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D2 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D3 = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D4 = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D5 = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D6 = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A2 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A6 = CLBLM_L_X12Y147_SLICE_X16Y147_B_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_AX = 1'b0;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B3 = CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B5 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B6 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_BX = CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C1 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C4 = CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C5 = CLBLM_L_X12Y147_SLICE_X17Y147_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_CX = CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D1 = CLBLM_L_X12Y147_SLICE_X17Y147_BQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D2 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D4 = CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_DX = CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A3 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A5 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_AX = 1'b0;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B2 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B3 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B5 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_BX = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C1 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C3 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C5 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_CX = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D1 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D3 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D5 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_DX = CLBLM_L_X12Y147_SLICE_X16Y147_BQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A1 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A2 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A3 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A4 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A5 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A6 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_AX = CLBLM_R_X15Y152_SLICE_X21Y152_CO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B1 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B2 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B3 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B4 = CLBLM_R_X15Y151_SLICE_X20Y151_BQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B5 = CLBLM_L_X16Y151_SLICE_X22Y151_C_XOR;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C3 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C4 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C5 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C6 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A4 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D1 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D2 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D3 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D4 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A6 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D6 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_AX = 1'b0;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B6 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A3 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_BX = 1'b0;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A4 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C6 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_AX = CLBLM_R_X15Y151_SLICE_X20Y151_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CIN = CLBLM_R_X11Y130_SLICE_X15Y130_COUT;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B2 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B3 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B4 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CX = 1'b0;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_BX = CLBLM_R_X15Y151_SLICE_X20Y151_CO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D6 = CLBLM_L_X12Y132_SLICE_X17Y132_A5Q;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C3 = CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C4 = CLBLM_L_X16Y153_SLICE_X22Y153_D_XOR;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_DX = 1'b0;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A6 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D2 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A2 = CLBLM_R_X3Y157_SLICE_X3Y157_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A3 = CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A4 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A5 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A6 = CLBLL_L_X2Y153_SLICE_X0Y153_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_AX = 1'b0;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_AX = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B6 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_BX = 1'b0;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_CE = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CIN = CLBLM_R_X11Y130_SLICE_X14Y130_COUT;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CX = 1'b0;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_DX = 1'b0;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A1 = CLBLL_L_X2Y153_SLICE_X0Y153_C5Q;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A2 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A3 = CLBLM_R_X3Y153_SLICE_X2Y153_CQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A4 = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A5 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_AX = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B1 = CLBLM_R_X3Y157_SLICE_X3Y157_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B2 = CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B3 = CLBLL_L_X2Y153_SLICE_X0Y153_D5Q;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B4 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B5 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B6 = CLBLM_R_X3Y153_SLICE_X2Y153_DQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_BX = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C1 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C3 = CLBLL_L_X2Y153_SLICE_X0Y153_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C4 = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C6 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_CE = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_CX = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D3 = CLBLL_L_X2Y153_SLICE_X0Y153_A5Q;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D4 = CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D5 = CLBLM_R_X3Y153_SLICE_X2Y153_BQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D6 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A2 = CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_DX = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A4 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A5 = CLBLM_L_X12Y147_SLICE_X17Y147_CQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A6 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_AX = CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B2 = CLBLM_L_X12Y147_SLICE_X17Y147_DQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B3 = CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B4 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B6 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_BX = CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C1 = CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C2 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C5 = CLBLM_L_X12Y148_SLICE_X17Y148_AQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_CIN = CLBLM_L_X12Y147_SLICE_X17Y147_COUT;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_CX = CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D2 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D3 = CLBLM_L_X12Y148_SLICE_X17Y148_BQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D5 = CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A1 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_DX = CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A2 = CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A4 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A5 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B2 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B4 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B5 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C1 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C2 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C4 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C5 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_CIN = CLBLM_L_X12Y147_SLICE_X16Y147_COUT;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D1 = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D2 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D4 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D6 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_A1 = CLBLM_L_X16Y150_SLICE_X22Y150_B_XOR;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_A2 = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_A3 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_A4 = CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_A5 = CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_A6 = CLBLM_R_X15Y150_SLICE_X21Y150_AO5;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_AX = CLBLM_R_X15Y152_SLICE_X21Y152_BO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_B1 = CLBLM_L_X16Y152_SLICE_X22Y152_B_XOR;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_B2 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_B3 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_B4 = CLBLM_R_X15Y152_SLICE_X21Y152_DO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_B5 = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_B6 = CLBLM_L_X16Y150_SLICE_X22Y150_A_XOR;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_BX = CLBLM_R_X15Y153_SLICE_X21Y153_CO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_C1 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_C2 = CLBLM_R_X15Y150_SLICE_X21Y150_AO5;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_C3 = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_C4 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D3 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_C5 = CLBLM_L_X16Y150_SLICE_X22Y150_B_XOR;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_C6 = CLBLM_L_X16Y152_SLICE_X22Y152_C_XOR;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D4 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D5 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_D1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_D2 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_D3 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_D4 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A6 = CLBLM_L_X12Y131_SLICE_X17Y131_A5Q;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_D5 = CLBLM_R_X15Y152_SLICE_X21Y152_AQ;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_AX = 1'b0;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_A1 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B6 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_A2 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_BX = 1'b0;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_A3 = CLBLM_R_X15Y152_SLICE_X20Y152_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C6 = CLBLM_L_X12Y132_SLICE_X17Y132_B5Q;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_AX = CLBLM_R_X15Y152_SLICE_X20Y152_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_CIN = CLBLM_R_X11Y131_SLICE_X15Y131_COUT;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_B1 = CLBLM_L_X16Y153_SLICE_X22Y153_B_XOR;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_B2 = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_B3 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_B4 = CLBLM_L_X16Y151_SLICE_X22Y151_A_XOR;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_B5 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_CX = 1'b0;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D6 = CLBLM_L_X12Y131_SLICE_X16Y131_A5Q;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_C3 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_C4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_DX = 1'b0;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_D1 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_D2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A2 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A3 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A6 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_D3 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_D4 = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A1 = CLBLM_R_X3Y157_SLICE_X3Y157_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A2 = CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A3 = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A4 = CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A5 = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_AX = 1'b0;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B1 = CLBLM_R_X3Y157_SLICE_X3Y157_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B4 = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B5 = CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B6 = CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B6 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CE = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CIN = CLBLM_R_X11Y131_SLICE_X14Y131_COUT;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CX = 1'b0;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D3 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_DX = 1'b0;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A1 = CLBLM_R_X3Y159_SLICE_X3Y159_CQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A2 = CLBLM_R_X3Y158_SLICE_X2Y158_A5Q;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A3 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A4 = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_AX = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B1 = CLBLM_R_X3Y155_SLICE_X2Y155_CQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B2 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B3 = CLBLM_R_X3Y154_SLICE_X2Y154_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B4 = CLBLM_R_X3Y155_SLICE_X2Y155_DQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B6 = CLBLM_R_X3Y155_SLICE_X2Y155_A5Q;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C1 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C2 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C3 = CLBLM_R_X3Y158_SLICE_X2Y158_CQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C4 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C5 = CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C6 = CLBLM_R_X3Y159_SLICE_X3Y159_CQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D1 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D2 = CLBLM_R_X3Y154_SLICE_X2Y154_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D3 = CLBLM_R_X3Y158_SLICE_X2Y158_A5Q;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D4 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D5 = CLBLM_R_X3Y155_SLICE_X2Y155_CQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D6 = CLBLM_R_X3Y155_SLICE_X2Y155_DQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A1 = CLBLM_L_X12Y148_SLICE_X17Y148_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A3 = CLBLM_L_X12Y149_SLICE_X16Y149_B_CY;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A6 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_AX = CLBLM_L_X12Y149_SLICE_X16Y149_B_CY;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B1 = CLBLM_L_X12Y148_SLICE_X17Y148_DQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B6 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X2Y139_SLICE_X1Y139_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_BX = 1'b0;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C1 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C2 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C5 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_CIN = CLBLM_L_X12Y148_SLICE_X17Y148_COUT;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_CX = 1'b0;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D1 = CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D2 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X2Y139_SLICE_X1Y139_BO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_DX = 1'b0;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A4 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_AX = 1'b0;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B3 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B6 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_BX = 1'b0;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C6 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_CIN = CLBLM_L_X12Y148_SLICE_X16Y148_COUT;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_CX = 1'b0;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D6 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_DX = 1'b0;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B2 = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLL_L_X2Y139_SLICE_X1Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A3 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A2 = CLBLM_R_X15Y152_SLICE_X21Y152_BQ;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A3 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A4 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A5 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B2 = CLBLM_L_X16Y150_SLICE_X22Y150_D_XOR;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B3 = CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B4 = CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B5 = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B6 = CLBLM_R_X15Y153_SLICE_X21Y153_AO5;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C2 = CLBLM_L_X16Y153_SLICE_X22Y153_A_XOR;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C3 = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C4 = CLBLM_R_X15Y153_SLICE_X21Y153_AO5;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C5 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C6 = CLBLM_L_X16Y150_SLICE_X22Y150_D_XOR;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D2 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D4 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_AX = 1'b0;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A2 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_BX = 1'b0;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C4 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_CIN = CLBLM_R_X11Y132_SLICE_X15Y132_COUT;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B1 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B4 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_CX = 1'b0;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D6 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_DX = 1'b0;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A2 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A5 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A6 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A1 = CLBLM_R_X3Y155_SLICE_X2Y155_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A2 = CLBLM_R_X3Y155_SLICE_X3Y155_BQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A3 = CLBLM_R_X3Y155_SLICE_X3Y155_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A4 = CLBLM_R_X3Y155_SLICE_X3Y155_CQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_AX = 1'b0;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_AX = CLBLM_R_X3Y159_SLICE_X3Y159_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B1 = CLBLM_R_X3Y159_SLICE_X3Y159_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B2 = CLBLM_R_X3Y155_SLICE_X3Y155_BQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B4 = CLBLM_R_X3Y155_SLICE_X3Y155_CQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B5 = CLBLM_R_X3Y155_SLICE_X2Y155_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B6 = CLBLM_L_X12Y132_SLICE_X17Y132_B5Q;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_BX = CLBLM_R_X3Y159_SLICE_X2Y159_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_BX = 1'b0;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C1 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C2 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C3 = CLBLM_R_X3Y155_SLICE_X2Y155_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C4 = CLBLM_R_X3Y159_SLICE_X3Y159_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C5 = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C6 = CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CIN = CLBLM_R_X11Y132_SLICE_X14Y132_COUT;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CX = 1'b0;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_CX = CLBLL_L_X2Y158_SLICE_X0Y158_CQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D2 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D3 = CLBLM_R_X3Y155_SLICE_X3Y155_DQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D4 = CLBLM_R_X3Y155_SLICE_X3Y155_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D5 = CLBLM_R_X3Y155_SLICE_X3Y155_BQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D6 = CLBLM_R_X3Y155_SLICE_X3Y155_CQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_DX = CLBLM_R_X3Y155_SLICE_X2Y155_AQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_DX = 1'b0;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A4 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A6 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_AX = CLBLM_R_X3Y158_SLICE_X2Y158_A5Q;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B1 = CLBLL_L_X2Y158_SLICE_X0Y158_CQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B2 = CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B5 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B6 = CLBLM_R_X3Y159_SLICE_X2Y159_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A1 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A2 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_BX = CLBLM_R_X3Y154_SLICE_X2Y154_AQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C1 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C2 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C3 = CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C4 = CLBLM_R_X3Y154_SLICE_X2Y154_AQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C5 = CLBLM_R_X3Y158_SLICE_X2Y158_A5Q;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C6 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A4 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_CX = CLBLM_R_X3Y159_SLICE_X3Y159_CQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D2 = CLBLM_R_X3Y155_SLICE_X2Y155_CQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D3 = CLBLM_R_X3Y155_SLICE_X2Y155_DQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D4 = CLBLM_R_X3Y155_SLICE_X2Y155_A5Q;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D5 = CLBLM_R_X3Y155_SLICE_X2Y155_BQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A1 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A4 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_DX = CLBLM_R_X3Y158_SLICE_X2Y158_CQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_AX = 1'b0;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B5 = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B1 = CLBLM_L_X12Y149_SLICE_X17Y149_DQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B5 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B6 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign RIOB33_X105Y125_IOB_X1Y125_O = CLBLM_L_X16Y133_SLICE_X22Y133_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_BX = 1'b0;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C1 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C5 = CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_CIN = CLBLM_L_X12Y149_SLICE_X17Y149_COUT;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_CX = 1'b0;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_DX = 1'b0;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A3 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A4 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A6 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B2 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B4 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B5 = CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B6 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C2 = CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C5 = CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C6 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D1 = CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D2 = CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D3 = CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D4 = CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D6 = CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A1 = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A2 = CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A3 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A4 = CLBLM_R_X11Y135_SLICE_X15Y135_CQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A5 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B1 = CLBLL_L_X26Y133_SLICE_X38Y133_DO5;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B2 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B3 = CLBLL_L_X26Y133_SLICE_X38Y133_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B4 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B6 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C1 = CLBLM_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C2 = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C3 = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C4 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C6 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D1 = CLBLM_R_X3Y126_SLICE_X2Y126_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D2 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D4 = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D5 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D6 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A2 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A3 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A4 = CLBLL_L_X26Y133_SLICE_X38Y133_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A5 = CLBLL_L_X26Y133_SLICE_X38Y133_CO5;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A6 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A1 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A2 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A4 = CLBLM_R_X3Y156_SLICE_X3Y156_BO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A5 = CLBLM_R_X3Y158_SLICE_X2Y158_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A6 = CLBLM_R_X3Y156_SLICE_X2Y156_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_AX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B1 = CLBLL_L_X26Y133_SLICE_X38Y133_BO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_AX = CLBLM_R_X3Y158_SLICE_X2Y158_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B2 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B1 = CLBLM_R_X3Y156_SLICE_X3Y156_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B2 = CLBLL_L_X2Y155_SLICE_X1Y155_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B3 = CLBLM_R_X3Y156_SLICE_X3Y156_CQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B5 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B6 = CLBLM_R_X3Y156_SLICE_X2Y156_CQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B6 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_BX = CLBLL_L_X2Y155_SLICE_X1Y155_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_BX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C1 = CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C2 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C3 = CLBLL_L_X2Y155_SLICE_X1Y155_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C4 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C5 = CLBLM_R_X3Y156_SLICE_X3Y156_DO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C6 = CLBLM_R_X3Y156_SLICE_X2Y156_BQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C5 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CE = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D1 = CLBLL_L_X26Y133_SLICE_X38Y133_CO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_CX = CLBLM_R_X3Y156_SLICE_X2Y156_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D1 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D2 = CLBLM_R_X3Y156_SLICE_X3Y156_CQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D3 = CLBLM_R_X3Y156_SLICE_X3Y156_BQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D4 = CLBLM_R_X3Y156_SLICE_X2Y156_CQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D5 = CLBLM_R_X3Y156_SLICE_X3Y156_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D6 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D4 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A1 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A3 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A4 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A5 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A6 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_AX = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B1 = CLBLM_R_X3Y159_SLICE_X2Y159_CQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B2 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B3 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B5 = CLBLM_R_X3Y158_SLICE_X2Y158_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B6 = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_BX = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C1 = CLBLM_R_X3Y156_SLICE_X3Y156_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C2 = CLBLM_R_X3Y156_SLICE_X2Y156_CQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C3 = CLBLL_L_X2Y155_SLICE_X1Y155_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C6 = CLBLM_R_X3Y156_SLICE_X2Y156_BQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_CX = CLBLM_R_X3Y159_SLICE_X2Y159_CQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D1 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D2 = CLBLM_R_X3Y158_SLICE_X2Y158_BQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D3 = CLBLM_R_X3Y158_SLICE_X2Y158_DQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D6 = CLBLM_R_X3Y157_SLICE_X2Y157_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A2 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A3 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A5 = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A6 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_AX = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B2 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B3 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B5 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B6 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_BX = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C1 = CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C2 = CLBLM_R_X15Y152_SLICE_X21Y152_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C3 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C5 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C6 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLL_L_X2Y147_SLICE_X0Y147_A5Q;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_CX = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D1 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D2 = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D4 = CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D6 = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A3 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A4 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A5 = CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A6 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B1 = CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B2 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B3 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B4 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B5 = CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B6 = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C1 = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C2 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C3 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C4 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C5 = CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C6 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A1 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A3 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A4 = CLBLM_L_X12Y131_SLICE_X16Y131_A5Q;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A5 = CLBLM_L_X12Y137_SLICE_X16Y137_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B1 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B2 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B3 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B5 = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B6 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C2 = CLBLM_R_X11Y135_SLICE_X15Y135_CQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C3 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C4 = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C5 = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C6 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D1 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D2 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D3 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D4 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D5 = CLBLM_R_X11Y135_SLICE_X15Y135_CQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A2 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A3 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A4 = CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A5 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A6 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A1 = CLBLM_R_X3Y157_SLICE_X2Y157_DQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A2 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A3 = CLBLM_R_X3Y157_SLICE_X3Y157_CQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A4 = CLBLM_R_X3Y157_SLICE_X2Y157_BQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A6 = CLBLM_R_X3Y157_SLICE_X2Y157_CQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B1 = CLBLL_L_X26Y133_SLICE_X38Y133_AO5;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_AX = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B1 = CLBLM_R_X3Y158_SLICE_X3Y158_DO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B2 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B3 = CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B4 = CLBLM_R_X3Y159_SLICE_X3Y159_BQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B5 = CLBLM_R_X3Y157_SLICE_X2Y157_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B6 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B6 = CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_BX = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C1 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C2 = CLBLM_R_X3Y157_SLICE_X3Y157_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C3 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C4 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C5 = CLBLM_R_X3Y157_SLICE_X3Y157_DO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C6 = CLBLM_R_X3Y157_SLICE_X2Y157_BQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C5 = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D1 = CLBLM_R_X11Y135_SLICE_X15Y135_CQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D2 = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_CX = CLBLM_R_X3Y157_SLICE_X3Y157_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D3 = CLBLM_R_X13Y135_SLICE_X18Y135_AO5;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D1 = CLBLM_R_X3Y157_SLICE_X2Y157_CQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D2 = CLBLM_R_X3Y157_SLICE_X3Y157_CQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D3 = CLBLM_R_X3Y157_SLICE_X3Y157_DQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D6 = CLBLM_R_X3Y157_SLICE_X2Y157_DQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D4 = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D5 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_DX = CLBLM_R_X3Y157_SLICE_X2Y157_BQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A1 = CLBLM_R_X3Y157_SLICE_X3Y157_AQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A2 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A3 = CLBLM_R_X3Y157_SLICE_X3Y157_AO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A4 = CLBLM_R_X3Y158_SLICE_X2Y158_BQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A5 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A6 = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_AX = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B1 = CLBLM_R_X3Y157_SLICE_X2Y157_BQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B2 = CLBLM_R_X3Y157_SLICE_X2Y157_DQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B4 = CLBLM_R_X3Y157_SLICE_X2Y157_CQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B5 = CLBLM_R_X3Y157_SLICE_X3Y157_AQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_BX = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C2 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C3 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_CX = CLBLM_R_X3Y158_SLICE_X2Y158_BQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D1 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D2 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D3 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D4 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D5 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D6 = 1'b1;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_DX = CLBLM_R_X3Y158_SLICE_X2Y158_DQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A2 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A3 = CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A4 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A5 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_AX = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B2 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B5 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C1 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C2 = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C4 = CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C5 = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C6 = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D3 = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D4 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D6 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A1 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A2 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A3 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A4 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B1 = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B2 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B3 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B4 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B5 = CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C2 = CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C3 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C5 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C6 = CLBLM_R_X13Y135_SLICE_X18Y135_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D1 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D3 = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A1 = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A2 = CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A3 = CLBLM_R_X13Y136_SLICE_X18Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A4 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A6 = CLBLM_R_X7Y136_SLICE_X9Y136_AO5;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A2 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A3 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A4 = CLBLM_R_X3Y159_SLICE_X2Y159_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A5 = CLBLM_R_X3Y158_SLICE_X3Y158_BO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A6 = CLBLM_R_X3Y159_SLICE_X3Y159_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B2 = CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B3 = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_AX = CLBLM_R_X3Y159_SLICE_X3Y159_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B2 = CLBLM_R_X3Y158_SLICE_X3Y158_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B3 = CLBLM_R_X3Y158_SLICE_X3Y158_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B5 = CLBLM_R_X3Y157_SLICE_X2Y157_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B6 = CLBLM_R_X3Y158_SLICE_X3Y158_CQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B6 = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_BX = CLBLM_R_X3Y159_SLICE_X2Y159_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C1 = CLBLM_R_X3Y157_SLICE_X2Y157_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C2 = CLBLM_R_X3Y158_SLICE_X3Y158_CQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C3 = CLBLM_R_X3Y158_SLICE_X3Y158_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C4 = CLBLM_R_X3Y159_SLICE_X3Y159_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C5 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_CE = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D1 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_CX = CLBLM_R_X3Y159_SLICE_X2Y159_DQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D2 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D1 = CLBLM_R_X3Y158_SLICE_X3Y158_CQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D2 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D3 = CLBLM_R_X3Y158_SLICE_X3Y158_DQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D4 = CLBLM_R_X3Y158_SLICE_X3Y158_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D5 = CLBLM_R_X3Y158_SLICE_X3Y158_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D6 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D4 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_DX = CLBLM_R_X3Y157_SLICE_X2Y157_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A6 = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_AX = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B2 = CLBLM_R_X3Y159_SLICE_X2Y159_DQ;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B3 = CLBLM_R_X3Y158_SLICE_X3Y158_CO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B4 = CLBLM_R_X3Y159_SLICE_X2Y159_BQ;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B5 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_BX = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C6 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_CX = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D6 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_DX = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A2 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A3 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A4 = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A5 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B1 = CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B2 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B3 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B4 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B5 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C1 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C4 = CLBLM_R_X7Y138_SLICE_X9Y138_AO5;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C5 = CLBLL_L_X26Y133_SLICE_X38Y133_BO5;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C6 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D1 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D2 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D3 = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D4 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D5 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C3 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A2 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A3 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A4 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A5 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A6 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C4 = CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C5 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B1 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B2 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B3 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B4 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B5 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B6 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C3 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C4 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C6 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D2 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D3 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D4 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A1 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A2 = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A3 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A4 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A5 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B1 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B2 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B3 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B4 = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B5 = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B6 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C5 = CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_CE = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D2 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A1 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A2 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A3 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A4 = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A5 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A6 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_A1 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_A2 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_A3 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_A4 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_A5 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_A6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_AX = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B1 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_AX = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B2 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_B1 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_B2 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_B3 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_B4 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_B5 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_B6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B6 = CLBLM_L_X16Y134_SLICE_X22Y134_CO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B1 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_BX = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_C1 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_C2 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_C3 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B2 = CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_C4 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_C5 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_C6 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B3 = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_CX = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D2 = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_CX = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D3 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_D1 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_D2 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_D3 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_D4 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_D5 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_D6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D4 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D5 = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_R_X3Y159_SLICE_X3Y159_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B6 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_A1 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_A2 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_A3 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_A4 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_A5 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_A6 = 1'b1;
  assign LIOB33_X0Y51_IOB_X0Y51_O = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign LIOB33_X0Y51_IOB_X0Y52_O = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_AX = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_B1 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_B2 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_B3 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_B4 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_B5 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_B6 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_BX = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_C1 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_C2 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_C3 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C2 = CLBLM_L_X10Y140_SLICE_X12Y140_AO5;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_C4 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_C5 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_C6 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C3 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C4 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_CX = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_D1 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_D2 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_D3 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_D4 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_D5 = 1'b1;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_D6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C6 = CLBLM_R_X13Y140_SLICE_X19Y140_BO6;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_DX = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_R_X3Y159_SLICE_X2Y159_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A1 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A3 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A4 = CLBLM_L_X16Y136_SLICE_X22Y136_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A6 = CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B1 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B3 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B4 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B6 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C1 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C2 = CLBLM_R_X5Y138_SLICE_X7Y138_CO5;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C3 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C4 = CLBLL_L_X26Y133_SLICE_X38Y133_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C5 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C6 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D5 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D1 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D3 = CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A1 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A2 = CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A3 = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A4 = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A5 = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A6 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_AX = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B1 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B2 = CLBLM_R_X13Y136_SLICE_X19Y136_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B3 = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B4 = CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B5 = CLBLM_R_X13Y133_SLICE_X19Y133_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B6 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_BX = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C1 = CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C2 = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C3 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C4 = CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C5 = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C6 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D6 = CLBLM_R_X13Y146_SLICE_X18Y146_C_XOR;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_CX = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D1 = CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D2 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D3 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D4 = CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D5 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D6 = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A1 = CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A3 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A4 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A5 = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A6 = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B1 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B2 = CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B3 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B4 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B5 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B6 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C2 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C3 = CLBLM_R_X13Y138_SLICE_X18Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C4 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C5 = CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D3 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D4 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D5 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D6 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_BI = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_CE = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_DI = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A2 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A3 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A4 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A5 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A6 = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B1 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B3 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B4 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B6 = CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C1 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C5 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D2 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D3 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D4 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D5 = CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D6 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A1 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A2 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A3 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A5 = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A6 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_B6 = CLBLM_R_X15Y152_SLICE_X20Y152_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B2 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B3 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B5 = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B6 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C1 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C2 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C3 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C4 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D2 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D4 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D5 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D6 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A1 = CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A2 = CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A3 = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A4 = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A5 = CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B1 = CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B3 = CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B4 = CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B5 = CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B6 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C3 = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C5 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_CE = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D2 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D4 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_BI = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CE = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_DI = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A1 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A2 = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A3 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A4 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A5 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B1 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B3 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B4 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B5 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C2 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C4 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C5 = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C6 = CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X2Y144_SLICE_X0Y144_A5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D2 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D3 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D5 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A1 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A2 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A3 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A5 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A6 = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B1 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B2 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B3 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B5 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B6 = CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C2 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C3 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C4 = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C5 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = CLBLM_L_X16Y133_SLICE_X22Y133_CQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_AO5;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D3 = CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D4 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D6 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = CLBLM_L_X16Y133_SLICE_X23Y133_DQ;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A1 = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A2 = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A3 = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A4 = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A6 = CLBLM_L_X12Y142_SLICE_X16Y142_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B1 = CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B3 = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B4 = CLBLM_R_X13Y140_SLICE_X18Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B5 = CLBLM_L_X12Y141_SLICE_X16Y141_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B6 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C1 = CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C2 = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C3 = CLBLM_R_X13Y140_SLICE_X18Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C4 = CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C5 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C6 = CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_CE = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D1 = CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D2 = CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D3 = CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D5 = CLBLM_R_X13Y140_SLICE_X18Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_AI = CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_BI = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CE = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CI = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_DI = 1'b0;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A1 = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A3 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A4 = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A5 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B1 = CLBLM_L_X12Y137_SLICE_X16Y137_CO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B2 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B3 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B5 = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C1 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C3 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C4 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C5 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C6 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D2 = CLBLM_L_X16Y137_SLICE_X22Y137_AO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D3 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D4 = CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D6 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A1 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A2 = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A3 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A4 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A5 = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A6 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B2 = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B5 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B6 = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C1 = CLBLL_L_X4Y136_SLICE_X5Y136_AO5;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C2 = CLBLM_L_X16Y137_SLICE_X23Y137_AO5;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C4 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C5 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C6 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D2 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D3 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D4 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D6 = CLBLM_R_X5Y137_SLICE_X7Y137_AO5;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A1 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A2 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A3 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A4 = CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A5 = CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_AX = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B1 = CLBLM_R_X11Y143_SLICE_X15Y143_A5Q;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B2 = CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B3 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B4 = CLBLM_R_X11Y141_SLICE_X15Y141_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B5 = CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_BX = CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C1 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C2 = CLBLM_R_X11Y140_SLICE_X15Y140_DQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C3 = CLBLM_R_X11Y141_SLICE_X15Y141_DQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C4 = CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_CX = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D1 = CLBLM_L_X12Y141_SLICE_X17Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D2 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D3 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D5 = CLBLM_R_X11Y141_SLICE_X15Y141_BO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_DX = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_AI = CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_BI = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_CE = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_CI = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_DI = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A1 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A2 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A4 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A5 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B6 = CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C2 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C5 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D3 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D5 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D6 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A2 = CLBLM_R_X15Y142_SLICE_X20Y142_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A3 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A5 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B2 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B3 = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B4 = CLBLM_R_X15Y140_SLICE_X21Y140_AO5;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C1 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C3 = CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C4 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C6 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D1 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D6 = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B6 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X2Y147_SLICE_X0Y147_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A1 = CLBLM_R_X11Y141_SLICE_X15Y141_DQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A2 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A3 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A4 = CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A5 = CLBLM_R_X11Y141_SLICE_X15Y141_CQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A6 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_AX = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B1 = CLBLM_R_X11Y140_SLICE_X15Y140_DQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B2 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B3 = CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B4 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B6 = CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C3 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_L_X2Y145_SLICE_X0Y145_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_BX = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C1 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C2 = CLBLM_R_X11Y143_SLICE_X15Y143_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C3 = CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C4 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C6 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C6 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_CX = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D1 = CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D3 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D4 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D6 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_DX = CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A4 = CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A5 = CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_AI = CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_BI = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = CLBLM_R_X13Y138_SLICE_X19Y138_CQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_CE = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_CI = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_DI = 1'b0;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = CLBLM_L_X16Y136_SLICE_X23Y136_DQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B5 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C1 = CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C2 = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A1 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A2 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A3 = CLBLL_L_X2Y131_SLICE_X0Y131_AQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A4 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A5 = CLBLL_L_X2Y131_SLICE_X0Y131_BQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A6 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_AX = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B1 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B2 = CLBLL_L_X2Y131_SLICE_X0Y131_BQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B5 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B6 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_BX = CLBLL_L_X4Y133_SLICE_X5Y133_F7AMUX_O;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C1 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C2 = CLBLL_L_X2Y131_SLICE_X0Y131_AQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C5 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C6 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_CE = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_BX = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A1 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A2 = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A3 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A4 = CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B2 = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B4 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B5 = CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B6 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C1 = CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C2 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C4 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C5 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C6 = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_CE = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_AX = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D2 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D3 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D4 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D5 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_CE = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A1 = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_AX = CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A3 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B2 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B5 = CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B6 = CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C1 = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C2 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C3 = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C4 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C5 = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C6 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D1 = CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D3 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D4 = CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D5 = CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A2 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A3 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A4 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_AX = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B1 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B2 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B3 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B4 = CLBLM_R_X11Y142_SLICE_X15Y142_F7BMUX_O;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C5 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B5 = CLBLM_R_X11Y142_SLICE_X15Y142_F7AMUX_O;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B6 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C1 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C3 = CLBLM_R_X11Y141_SLICE_X15Y141_DQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C4 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C5 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C6 = CLBLM_R_X11Y136_SLICE_X14Y136_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_A2 = CLBLM_L_X16Y133_SLICE_X22Y133_AQ;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_A3 = CLBLM_L_X16Y133_SLICE_X23Y133_AQ;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_A6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D2 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_B1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_B2 = CLBLM_L_X16Y133_SLICE_X22Y133_BQ;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_B4 = CLBLM_L_X16Y133_SLICE_X23Y133_BQ;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_B6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A1 = CLBLM_R_X15Y141_SLICE_X20Y141_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A2 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_C1 = CLBLM_L_X16Y134_SLICE_X23Y134_AQ;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_C4 = CLBLM_L_X16Y133_SLICE_X23Y133_CQ;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_C5 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_C6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A4 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A5 = CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B1 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B2 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B3 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B4 = CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_D1 = CLBLM_L_X16Y133_SLICE_X22Y133_CQ;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_D3 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_D5 = CLBLM_L_X16Y133_SLICE_X23Y133_DQ;
  assign CLBLL_L_X26Y133_SLICE_X38Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C1 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C2 = CLBLM_L_X10Y137_SLICE_X13Y137_CQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C3 = CLBLM_R_X11Y140_SLICE_X15Y140_DQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C4 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C5 = CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C6 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D1 = CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D2 = CLBLM_R_X11Y143_SLICE_X15Y143_A5Q;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D3 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D4 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D6 = CLBLM_L_X10Y137_SLICE_X13Y137_BQ;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_A1 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_A2 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_A3 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_A4 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_A5 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_A6 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_B1 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_B2 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_B3 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_B4 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_B5 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_B6 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_C1 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_C2 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_C3 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_C4 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_C5 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_C6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A6 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_D1 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_D2 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_D3 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_D4 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_D5 = 1'b1;
  assign CLBLL_L_X26Y133_SLICE_X39Y133_D6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A1 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A2 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B2 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B4 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B5 = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C3 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C5 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C6 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_AX = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C2 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D2 = CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C3 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D5 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_CE = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A1 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A2 = CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B2 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B4 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B6 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C2 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C3 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D2 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D4 = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D6 = 1'b1;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A6 = 1'b1;
  assign LIOI3_SING_X0Y50_OLOGIC_X0Y50_T1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A2 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B1 = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B2 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B3 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B5 = CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B6 = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C2 = CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C3 = CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C4 = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C5 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C6 = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X2Y143_SLICE_X0Y143_AQ;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A2 = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A3 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A4 = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A5 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_AX = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B1 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B4 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B5 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B6 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C1 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C2 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_AX = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C3 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C4 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C5 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D2 = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_CE = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A3 = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_AX = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B1 = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B5 = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C2 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C3 = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C4 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C6 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D3 = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D5 = CLBLL_L_X4Y141_SLICE_X5Y141_DQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D6 = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_D = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_D = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A1 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A5 = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B1 = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B2 = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B3 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B4 = CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B6 = CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C2 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C3 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_A2 = CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_A5 = CLBLM_L_X16Y135_SLICE_X23Y135_AQ;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_A6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C4 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C6 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_B1 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_B2 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_B3 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_B4 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_B5 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_B6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D2 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_C1 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_C2 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_C3 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_C4 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_C5 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_C6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A1 = CLBLM_L_X12Y147_SLICE_X16Y147_BQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A2 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A4 = CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A5 = CLBLM_L_X12Y144_SLICE_X16Y144_BO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A6 = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_D1 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_D2 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_D3 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_D4 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_D5 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X38Y135_D6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B1 = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B2 = CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B3 = CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B4 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B6 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C1 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C3 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C6 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D1 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D2 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D3 = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D4 = CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D6 = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_A1 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_A2 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_A3 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_A4 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_A5 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_A6 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_B1 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_B2 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_B3 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_B4 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_B5 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_B6 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_C1 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_C2 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_C3 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_C4 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_C5 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_C6 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_D1 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_D2 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_D3 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_D4 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_D5 = 1'b1;
  assign CLBLL_L_X26Y135_SLICE_X39Y135_D6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C5 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A2 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A3 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A4 = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A6 = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_AX = CLBLM_R_X15Y141_SLICE_X20Y141_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B1 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B5 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B6 = CLBLM_L_X8Y142_SLICE_X11Y142_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_BX = CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C1 = CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C3 = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C5 = CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C6 = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D2 = CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D3 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D4 = CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D5 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D6 = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A1 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A2 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A4 = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A5 = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A6 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B1 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B2 = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B5 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B6 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C1 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C2 = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C3 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C5 = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C6 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D1 = CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D2 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D3 = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D4 = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D6 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A1 = CLBLM_R_X13Y147_SLICE_X19Y147_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A2 = CLBLM_R_X13Y148_SLICE_X18Y148_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A4 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A5 = CLBLM_R_X13Y146_SLICE_X19Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A6 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B1 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B2 = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B3 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B4 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B5 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B6 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A2 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A3 = CLBLM_L_X16Y136_SLICE_X23Y136_DQ;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A4 = CLBLM_L_X16Y139_SLICE_X22Y139_BQ;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C2 = CLBLM_R_X13Y146_SLICE_X18Y146_D_XOR;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B2 = CLBLM_L_X16Y136_SLICE_X23Y136_CQ;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B5 = CLBLM_L_X16Y136_SLICE_X23Y136_BQ;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C6 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D3 = CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D4 = CLBLM_R_X13Y146_SLICE_X18Y146_A_XOR;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A1 = CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A2 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A3 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A4 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A5 = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A6 = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B1 = CLBLM_R_X15Y149_SLICE_X20Y149_AO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B2 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B4 = CLBLM_L_X12Y144_SLICE_X16Y144_BO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B6 = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C2 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C4 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C5 = CLBLM_R_X13Y146_SLICE_X18Y146_B_XOR;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C6 = CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D2 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D5 = CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B6 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B3 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_A6 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_B6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_C6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X0Y135_D6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A1 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A1 = CLBLM_R_X5Y141_SLICE_X7Y141_CQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A4 = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A5 = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A6 = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A4 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_A6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B3 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B5 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B6 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C1 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C2 = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C3 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C4 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C6 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C2 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_C6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_CE = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D1 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D2 = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D3 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D1 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D4 = CLBLL_L_X4Y141_SLICE_X5Y141_DQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D5 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D6 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D5 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_D6 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A2 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A4 = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A5 = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A6 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B1 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B2 = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B4 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B5 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C2 = CLBLM_R_X13Y146_SLICE_X19Y146_AO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C1 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C2 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C3 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C5 = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C6 = CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C4 = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C5 = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D2 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D3 = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D4 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D5 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D6 = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B6 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A1 = CLBLM_L_X12Y147_SLICE_X16Y147_CQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A2 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A3 = CLBLM_R_X13Y146_SLICE_X19Y146_AO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A4 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A5 = CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A6 = CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_AX = CLBLM_L_X12Y147_SLICE_X16Y147_DQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B2 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B4 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B5 = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C1 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D4 = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C1 = CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C2 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C2 = CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C4 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C5 = CLBLM_R_X13Y146_SLICE_X19Y146_AO5;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C3 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C6 = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D5 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D6 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D1 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C5 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D4 = CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D6 = CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A1 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A2 = CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A3 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A4 = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A5 = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A6 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_C1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B3 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B4 = CLBLM_R_X13Y147_SLICE_X18Y147_A_XOR;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B6 = CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C1 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C2 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C3 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C4 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C5 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C6 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_C2 = CLBLM_R_X15Y152_SLICE_X20Y152_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D2 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D3 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D5 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B1 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B3 = CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_D = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_D = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B6 = CLBLM_L_X10Y137_SLICE_X13Y137_DQ;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLL_L_X2Y147_SLICE_X0Y147_A5Q;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C5 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C6 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C1 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A1 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A2 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A3 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A4 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A5 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C3 = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B1 = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B2 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B3 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B4 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B5 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B6 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A4 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C6 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C1 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C2 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C3 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C4 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C5 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C6 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A1 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A2 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A3 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A4 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A5 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A6 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_AX = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B2 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B3 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C6 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D2 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D3 = CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D4 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D5 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D6 = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A1 = CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A2 = CLBLM_R_X13Y146_SLICE_X19Y146_AO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A3 = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A4 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A5 = CLBLM_L_X12Y147_SLICE_X16Y147_DQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A6 = CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_A2 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_A3 = CLBLM_L_X16Y139_SLICE_X22Y139_AQ;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_A4 = CLBLM_L_X16Y138_SLICE_X23Y138_AQ;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_A6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D6 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_AX = CLBLM_L_X12Y147_SLICE_X16Y147_CQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B1 = CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_B1 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_B2 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_B3 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_B4 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_B5 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_B6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B6 = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C1 = CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_C1 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_C2 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_C3 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_C4 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_C5 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C6 = CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D2 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A2 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A6 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_D3 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_D5 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_D6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_AX = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B2 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X38Y138_D4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B6 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_BX = 1'b0;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C3 = CLBLL_L_X26Y133_SLICE_X38Y133_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C6 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B1 = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B2 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B3 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B5 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_CX = 1'b0;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D3 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_A1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D6 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_A2 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_A3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_DX = 1'b0;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_A4 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_A5 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_A6 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_B1 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_B2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A3 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A5 = CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A6 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_B3 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_B4 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_B5 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_B6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B1 = CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B2 = CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B3 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B5 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B6 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_C1 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_C2 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_C6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C1 = CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C2 = CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C3 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C6 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_D4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CE = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A2 = CLBLL_L_X2Y137_SLICE_X0Y137_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A3 = CLBLL_L_X2Y137_SLICE_X0Y137_AQ;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A4 = CLBLL_L_X2Y138_SLICE_X0Y138_C_XOR;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A5 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A6 = 1'b1;
  assign CLBLL_L_X26Y138_SLICE_X39Y138_D5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D6 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B4 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B5 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_BX = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C1 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C2 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C3 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C4 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C5 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_C6 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_CE = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D1 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D2 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D3 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D4 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D5 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_D6 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A1 = CLBLL_L_X2Y139_SLICE_X0Y139_A_XOR;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A2 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A3 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A4 = CLBLL_L_X2Y138_SLICE_X0Y138_D_XOR;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A5 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_A6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A1 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B1 = CLBLM_R_X3Y137_SLICE_X3Y137_DQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A3 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B2 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A4 = CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A5 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B3 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B4 = CLBLL_L_X2Y139_SLICE_X0Y139_B_XOR;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B5 = CLBLL_L_X2Y139_SLICE_X0Y139_C_XOR;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_B6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B3 = CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B4 = CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B5 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B6 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C1 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C2 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C3 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C4 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C5 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_C6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C1 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C3 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C4 = CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C6 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D1 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D2 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D3 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D4 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D5 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X1Y137_D6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D1 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D2 = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D3 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D4 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D5 = CLBLM_R_X3Y141_SLICE_X3Y141_DQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D6 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A1 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A2 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A4 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A5 = CLBLM_R_X5Y141_SLICE_X7Y141_CQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B1 = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B2 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B3 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B4 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B5 = CLBLM_R_X5Y141_SLICE_X7Y141_CQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B6 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C1 = CLBLM_R_X5Y141_SLICE_X7Y141_CQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C2 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C3 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C5 = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D1 = CLBLM_R_X5Y141_SLICE_X7Y141_CQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D2 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D3 = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D4 = CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_D = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A3 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A5 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B2 = CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B4 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B5 = CLBLM_R_X15Y150_SLICE_X20Y150_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B6 = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C1 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C6 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D1 = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D6 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D2 = CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D4 = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A6 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D6 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_AX = 1'b0;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A1 = CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B6 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A2 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A3 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_BX = 1'b0;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A4 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C6 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B3 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_CIN = CLBLM_R_X5Y128_SLICE_X7Y128_COUT;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B4 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B5 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C1 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_CX = 1'b0;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D6 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C4 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_DX = 1'b0;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C6 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D1 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A1 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A3 = CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A5 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A6 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D3 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D4 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B1 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B2 = CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B3 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B4 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B5 = CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B6 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A6 = CLBLL_L_X2Y140_SLICE_X1Y140_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C1 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_AX = 1'b0;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C2 = CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B2 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B3 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B5 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B6 = CLBLL_L_X2Y140_SLICE_X1Y140_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C3 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C4 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_BX = CLBLL_L_X2Y140_SLICE_X1Y140_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C6 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C6 = CLBLL_L_X2Y140_SLICE_X1Y140_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D1 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D2 = CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D3 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D4 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D5 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D6 = CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_CX = 1'b0;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D6 = CLBLL_L_X2Y140_SLICE_X1Y140_DQ;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_DX = 1'b0;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A1 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A2 = CLBLL_L_X2Y138_SLICE_X1Y138_BQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A3 = CLBLL_L_X2Y138_SLICE_X1Y138_AQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A4 = CLBLL_L_X2Y138_SLICE_X0Y138_A_XOR;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A5 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_AX = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A1 = CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A2 = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_BX = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A3 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_CE = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_AX = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B1 = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B2 = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B3 = CLBLM_R_X7Y145_SLICE_X8Y145_AO5;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B4 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C4 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C5 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C6 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D2 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D4 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D5 = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D6 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_D = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A1 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A3 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A4 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A5 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A6 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_AX = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A2 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A3 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A4 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A5 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B2 = CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B3 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B4 = CLBLM_R_X15Y151_SLICE_X20Y151_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B5 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign LIOI3_SING_X0Y199_ILOGIC_X0Y199_D = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C1 = CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C2 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C3 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C4 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C5 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C6 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D1 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D2 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D4 = CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A6 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D6 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_AX = 1'b0;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B6 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A2 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A3 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_BX = 1'b0;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A4 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C6 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CIN = CLBLM_R_X5Y129_SLICE_X7Y129_COUT;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B1 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B2 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B3 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B4 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B5 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CX = 1'b0;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D6 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C3 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C4 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_DX = 1'b0;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C6 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D2 = CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A3 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A4 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D4 = CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_AX = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D6 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A6 = CLBLL_L_X2Y141_SLICE_X1Y141_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_AX = 1'b0;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B6 = CLBLL_L_X2Y141_SLICE_X1Y141_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_BX = 1'b0;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_BX = 1'b0;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C6 = CLBLL_L_X2Y141_SLICE_X1Y141_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CX = 1'b0;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_CIN = CLBLL_L_X2Y138_SLICE_X0Y138_COUT;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D6 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_CX = 1'b0;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D6 = CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_DX = 1'b0;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_DX = 1'b0;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A1 = CLBLL_L_X2Y140_SLICE_X0Y140_B_XOR;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A2 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A3 = CLBLL_L_X2Y139_SLICE_X1Y139_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A4 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A5 = CLBLL_L_X2Y140_SLICE_X0Y140_C_XOR;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D3 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_AX = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B1 = CLBLL_L_X2Y141_SLICE_X0Y141_A_XOR;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B2 = CLBLL_L_X2Y139_SLICE_X1Y139_BQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B3 = CLBLL_L_X2Y140_SLICE_X0Y140_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B4 = CLBLL_L_X2Y140_SLICE_X0Y140_D_XOR;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B5 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B6 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_BX = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C1 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C2 = CLBLL_L_X2Y139_SLICE_X1Y139_CQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C3 = CLBLL_L_X2Y139_SLICE_X1Y139_DQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C4 = CLBLL_L_X2Y141_SLICE_X0Y141_C_XOR;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C5 = CLBLL_L_X2Y141_SLICE_X0Y141_B_XOR;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C6 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_CE = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A4 = CLBLM_R_X15Y143_SLICE_X20Y143_AO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A5 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A6 = CLBLM_L_X8Y149_SLICE_X11Y149_F7AMUX_O;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_CX = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D1 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D2 = CLBLL_L_X2Y140_SLICE_X0Y140_A_XOR;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D3 = CLBLL_L_X2Y139_SLICE_X0Y139_D_XOR;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D4 = CLBLL_L_X2Y140_SLICE_X0Y140_BQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D5 = CLBLL_L_X2Y140_SLICE_X0Y140_CQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D6 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B4 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_DX = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C1 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C2 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C4 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C6 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D1 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D2 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D4 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A4 = CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A5 = CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D6 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B1 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D1 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D2 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D4 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D6 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A4 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_A6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_AX = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_BX = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_CIN = CLBLM_R_X5Y130_SLICE_X7Y130_COUT;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_CX = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A6 = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_DX = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A6 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A1 = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A2 = CLBLL_L_X2Y142_SLICE_X1Y142_AQ;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_AX = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_AX = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B1 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B4 = CLBLL_L_X2Y142_SLICE_X1Y142_BQ;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_BX = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_BX = 1'b0;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C3 = CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C4 = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C6 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_CE = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_CIN = CLBLL_L_X2Y139_SLICE_X0Y139_COUT;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C6 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CIN = CLBLM_R_X5Y130_SLICE_X6Y130_COUT;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CX = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_CX = 1'b0;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D6 = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_DX = 1'b0;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D6 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_DX = 1'b0;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B6 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A2 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A3 = CLBLL_L_X2Y140_SLICE_X1Y140_AQ;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A4 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A5 = CLBLL_L_X4Y142_SLICE_X4Y142_F7AMUX_O;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A6 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_AX = 1'b0;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B1 = CLBLL_L_X2Y144_SLICE_X1Y144_AO5;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B2 = CLBLL_L_X2Y140_SLICE_X1Y140_BQ;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B3 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B4 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B5 = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B6 = CLBLL_L_X4Y141_SLICE_X4Y141_F7AMUX_O;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_BX = CLBLL_L_X2Y144_SLICE_X1Y144_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C1 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C2 = CLBLL_L_X2Y140_SLICE_X1Y140_CQ;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C4 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C5 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_CE = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A3 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_CX = 1'b0;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D2 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D3 = CLBLL_L_X2Y140_SLICE_X1Y140_DQ;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D4 = CLBLM_R_X5Y141_SLICE_X7Y141_F7AMUX_O;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D5 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_DX = 1'b0;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C3 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D3 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A3 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B3 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A6 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C3 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D3 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B4 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B6 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_BX = 1'b0;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_D = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_D = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A2 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A3 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A4 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A5 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A6 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B1 = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B2 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B4 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B5 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B6 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C1 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C2 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C3 = CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C4 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C5 = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CIN = CLBLM_R_X5Y131_SLICE_X6Y131_COUT;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C6 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C4 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D1 = CLBLM_R_X5Y131_SLICE_X7Y131_A_CY;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D2 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D3 = CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D6 = CLBLM_R_X5Y133_SLICE_X6Y133_D_CY;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOB33_X105Y123_IOB_X1Y124_O = CLBLM_L_X16Y133_SLICE_X23Y133_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A2 = CLBLL_L_X2Y141_SLICE_X1Y141_D_XOR;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A3 = CLBLL_L_X2Y143_SLICE_X1Y143_AQ;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_AX = 1'b0;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B6 = CLBLL_L_X2Y143_SLICE_X1Y143_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_AX = 1'b0;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_BX = 1'b0;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C6 = CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_CE = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_CIN = CLBLL_L_X2Y140_SLICE_X0Y140_COUT;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_CX = 1'b0;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C6 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CX = 1'b0;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_DX = 1'b0;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D4 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D6 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_DX = 1'b0;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B1 = CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B2 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A1 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A2 = CLBLM_R_X5Y143_SLICE_X7Y143_F7AMUX_O;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A3 = CLBLL_L_X2Y141_SLICE_X1Y141_AQ;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A4 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_AX = 1'b0;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B1 = CLBLM_R_X5Y142_SLICE_X7Y142_F7AMUX_O;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B2 = CLBLL_L_X2Y141_SLICE_X1Y141_BQ;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B3 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B4 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B5 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B6 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_BX = 1'b0;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C1 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C2 = CLBLM_R_X5Y141_SLICE_X6Y141_F7AMUX_O;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C4 = CLBLL_L_X2Y141_SLICE_X1Y141_CQ;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C5 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_CE = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_CIN = CLBLL_L_X2Y140_SLICE_X1Y140_COUT;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A3 = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_CX = 1'b0;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A5 = CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D1 = CLBLL_L_X2Y141_SLICE_X0Y141_AQ;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D2 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D3 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D4 = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D5 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D6 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_AX = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_DX = 1'b0;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C2 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C3 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C4 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C5 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D2 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D3 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D4 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D5 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A2 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B2 = CLBLM_L_X16Y142_SLICE_X22Y142_AO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B3 = CLBLM_R_X5Y151_SLICE_X6Y151_BO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B4 = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B5 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B6 = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C3 = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B6 = CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B2 = CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A6 = CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D6 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A2 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A3 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A4 = CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A5 = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_AX = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B2 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B3 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B3 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B4 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B5 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B6 = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B4 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C1 = CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C2 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B5 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C3 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C4 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C5 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C6 = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B6 = CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D1 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D2 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D3 = CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D4 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D5 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D6 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_AX = CLBLL_L_X2Y142_SLICE_X1Y142_D_XOR;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A6 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_AX = 1'b0;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_CE = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C4 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_BX = 1'b0;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C6 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_CE = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_CIN = CLBLM_R_X5Y132_SLICE_X6Y132_COUT;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_CX = 1'b0;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_DX = 1'b0;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A2 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A3 = CLBLL_L_X2Y142_SLICE_X1Y142_AQ;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A4 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A5 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A6 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D6 = CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_AX = 1'b0;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B1 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B2 = CLBLL_L_X2Y142_SLICE_X1Y142_BQ;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B3 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B4 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B5 = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B6 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_BX = 1'b0;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C1 = CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C2 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C3 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C4 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_CE = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_CIN = CLBLL_L_X2Y141_SLICE_X1Y141_COUT;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D3 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_CX = 1'b0;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D1 = CLBLL_L_X2Y142_SLICE_X0Y142_AQ;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D2 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D3 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D4 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D5 = CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_DX = 1'b0;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A1 = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A2 = CLBLM_R_X5Y150_SLICE_X7Y150_CO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A4 = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A6 = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C4 = CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D6 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOB33_X105Y127_IOB_X1Y127_O = CLBLM_L_X16Y133_SLICE_X22Y133_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A1 = CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A2 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A3 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A4 = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A5 = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A6 = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B1 = CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B2 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B4 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C1 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C2 = CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C3 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C4 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C5 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C6 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D2 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A2 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D6 = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A1 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A2 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A3 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C6 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_CE = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B1 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B2 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B3 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B5 = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C3 = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C4 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D2 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D6 = 1'b1;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_D = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_D = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B4 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A1 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A2 = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A3 = CLBLL_L_X2Y143_SLICE_X1Y143_AQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A4 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A5 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A6 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_AX = 1'b0;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B1 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B2 = CLBLL_L_X2Y143_SLICE_X1Y143_BQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B3 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B4 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B5 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B6 = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D3 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_BX = 1'b0;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B5 = CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C1 = CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C2 = CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C4 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C5 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C6 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_CE = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_CIN = CLBLL_L_X2Y142_SLICE_X1Y142_COUT;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_CX = 1'b0;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D1 = CLBLL_L_X2Y142_SLICE_X1Y142_C_XOR;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_DX = 1'b0;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A4 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B4 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C4 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D4 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A1 = CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A4 = CLBLM_R_X5Y150_SLICE_X7Y150_CO5;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A6 = CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B1 = CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B6 = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D4 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOB33_X105Y129_IOB_X1Y130_O = CLBLM_L_X16Y134_SLICE_X23Y134_AQ;
  assign RIOB33_X105Y129_IOB_X1Y129_O = CLBLM_L_X16Y133_SLICE_X23Y133_CQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A1 = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A3 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A4 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A5 = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A6 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B1 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B2 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B3 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B4 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B5 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C3 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C3 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C5 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C6 = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D1 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D2 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A5 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_BX = CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A6 = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C6 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_CE = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B1 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B2 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B3 = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B4 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B5 = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C1 = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C5 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D3 = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D5 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A1 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A2 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A3 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A4 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A6 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B1 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B2 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B3 = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B5 = CLBLL_L_X2Y144_SLICE_X1Y144_AO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B6 = CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C1 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C2 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C4 = CLBLL_L_X2Y144_SLICE_X1Y144_AO5;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C5 = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C6 = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D6 = 1'b1;
  assign RIOB33_X105Y131_IOB_X1Y132_O = CLBLM_L_X16Y133_SLICE_X22Y133_CQ;
  assign RIOB33_X105Y131_IOB_X1Y131_O = CLBLM_L_X16Y133_SLICE_X23Y133_DQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A1 = CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A3 = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A5 = CLBLM_R_X5Y136_SLICE_X7Y136_DQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B1 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B2 = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B4 = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B5 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C2 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C3 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C5 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C6 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A1 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D3 = CLBLM_R_X5Y136_SLICE_X7Y136_DQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D4 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_CE = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A2 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A3 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A4 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A5 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B5 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C2 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C3 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C4 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C6 = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B1 = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B2 = CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D2 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D3 = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D4 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D5 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B3 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_A1 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_A2 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_A3 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_A4 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_A5 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_A6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A1 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A2 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A3 = CLBLL_L_X2Y144_SLICE_X1Y144_BO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A5 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A6 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_B1 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B6 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_B5 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_B6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C6 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_C6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_D1 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_D2 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_D3 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_D4 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X23Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D6 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_A1 = CLBLM_R_X15Y131_SLICE_X21Y131_CQ;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_A2 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_A3 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_A4 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_A5 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_A6 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_B1 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_B2 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_B3 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_B4 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_B5 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C5 = CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C6 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_C1 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_C2 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_C3 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_C4 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_C5 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_C6 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_CE = CLBLM_L_X12Y129_SLICE_X17Y129_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CE = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_D1 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_D2 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_D3 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_D4 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_D5 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_D6 = 1'b1;
  assign CLBLM_L_X16Y131_SLICE_X22Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_D = LIOB33_X0Y165_IOB_X0Y166_I;
  assign RIOB33_X105Y133_IOB_X1Y134_O = CLBLM_L_X16Y134_SLICE_X22Y134_BQ;
  assign RIOB33_X105Y133_IOB_X1Y133_O = CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_D = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B3 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B6 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A1 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A2 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A3 = LIOB33_X0Y183_IOB_X0Y184_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A5 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C3 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B1 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C4 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B2 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B3 = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B5 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C5 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C6 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C2 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C3 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C5 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D1 = CLBLM_R_X15Y140_SLICE_X21Y140_DO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D2 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D3 = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A4 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D5 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D6 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A5 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A1 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A2 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A4 = CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A5 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_AX = CLBLM_R_X15Y140_SLICE_X21Y140_DO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B2 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B3 = CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B6 = CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_BX = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C2 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C3 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C4 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C5 = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C6 = CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B2 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B3 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_CX = CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D3 = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D4 = CLBLM_R_X5Y137_SLICE_X6Y137_AO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D5 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D6 = CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C1 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C2 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign RIOB33_X105Y135_IOB_X1Y136_O = CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  assign RIOB33_X105Y135_IOB_X1Y135_O = CLBLM_L_X16Y135_SLICE_X23Y135_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C5 = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A4 = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A6 = CLBLM_R_X7Y145_SLICE_X8Y145_AO5;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B5 = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B6 = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A1 = CLBLM_R_X7Y138_SLICE_X8Y138_B_XOR;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A2 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A4 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A5 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_AX = CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B2 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B3 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B4 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B5 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_BX = CLBLM_R_X5Y138_SLICE_X7Y138_CO5;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A1 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C1 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C2 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C3 = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_CE = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A1 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A2 = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A3 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A4 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B1 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B2 = CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B3 = CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B4 = CLBLM_R_X15Y143_SLICE_X21Y143_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B5 = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B6 = CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C1 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C2 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C3 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C4 = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C5 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C6 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D2 = CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D3 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D4 = CLBLM_R_X15Y143_SLICE_X21Y143_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A6 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_A2 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_A3 = CLBLM_L_X16Y133_SLICE_X23Y133_AQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B6 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_A5 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C6 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_B5 = CLBLM_L_X16Y133_SLICE_X23Y133_BQ;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_C2 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_C3 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_C4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_C5 = CLBLM_L_X16Y133_SLICE_X23Y133_CQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D6 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_D3 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_D4 = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_D5 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_D6 = CLBLM_L_X16Y133_SLICE_X23Y133_DQ;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y133_SLICE_X23Y133_D2 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_A1 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_A2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_A3 = CLBLM_L_X16Y133_SLICE_X22Y133_AQ;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_A4 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign RIOB33_X105Y137_IOB_X1Y137_O = CLBLM_L_X16Y136_SLICE_X23Y136_BQ;
  assign RIOB33_X105Y137_IOB_X1Y138_O = CLBLM_L_X16Y136_SLICE_X23Y136_CQ;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_B2 = CLBLM_L_X16Y133_SLICE_X22Y133_BQ;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_B3 = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_B4 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_B5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_B6 = CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_C2 = CLBLM_L_X16Y133_SLICE_X22Y133_CQ;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_C3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_C4 = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_C5 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_C6 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_D1 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_D2 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_D3 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_D4 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_D5 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_D6 = 1'b1;
  assign CLBLM_L_X16Y133_SLICE_X22Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A2 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A3 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A6 = 1'b1;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_D = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_AX = CLBLM_R_X15Y142_SLICE_X20Y142_AO5;
  assign LIOI3_X0Y167_ILOGIC_X0Y167_D = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B1 = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B4 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B6 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_BX = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C1 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C3 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C4 = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C6 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D1 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D2 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D3 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D4 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D6 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A3 = CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A4 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A5 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B1 = CLBLL_L_X4Y141_SLICE_X5Y141_CQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B2 = CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B6 = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C2 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C3 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C4 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C5 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C6 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign LIOB33_X0Y53_IOB_X0Y53_O = CLBLL_L_X4Y135_SLICE_X5Y135_B5Q;
  assign LIOB33_X0Y53_IOB_X0Y54_O = CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A4 = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D1 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D2 = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B3 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B4 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_A2 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_A3 = CLBLM_L_X16Y134_SLICE_X23Y134_AQ;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_A4 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C3 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C6 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_B1 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_B4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_B5 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_B6 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_C1 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_C6 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D6 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_D1 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_D2 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_D3 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_D4 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_D5 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_D6 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X23Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_A2 = CLBLM_L_X16Y134_SLICE_X22Y134_BQ;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_A4 = CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_A6 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_B1 = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_B2 = CLBLM_L_X16Y134_SLICE_X22Y134_BQ;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_B4 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_B5 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_C1 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_C2 = CLBLM_L_X16Y134_SLICE_X22Y134_AO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_C3 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_C4 = CLBLM_L_X16Y134_SLICE_X22Y134_AO5;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_C6 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_D1 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_D2 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_D3 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_D4 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_D5 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_D6 = 1'b1;
  assign CLBLM_L_X16Y134_SLICE_X22Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A1 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A2 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A3 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A5 = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A6 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B4 = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C1 = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C2 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D1 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D2 = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D3 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D4 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D5 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D6 = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A1 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A3 = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A4 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A6 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B2 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B3 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B4 = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B6 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B3 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C1 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C3 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C6 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_CE = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A1 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A2 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A4 = CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A6 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A1 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A2 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A3 = CLBLM_L_X16Y135_SLICE_X23Y135_AQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B1 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B2 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B3 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_B5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C1 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C2 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C3 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_C6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D1 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D2 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D3 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_D6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X23Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A3 = CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A4 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A5 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_A6 = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B2 = CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B4 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B5 = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_B6 = CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C1 = CLBLM_L_X16Y136_SLICE_X22Y136_BQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C2 = CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C3 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_C6 = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D1 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D2 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D3 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D4 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D5 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_D6 = 1'b1;
  assign CLBLM_L_X16Y135_SLICE_X22Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D5 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C6 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A1 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A2 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A3 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A5 = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A6 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_AX = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B1 = CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B2 = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B3 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B5 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B6 = CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  assign LIOB33_X0Y57_IOB_X0Y57_O = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign LIOB33_X0Y57_IOB_X0Y58_O = CLBLM_R_X5Y136_SLICE_X7Y136_DQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C1 = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C5 = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C6 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_CE = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D1 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D2 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D3 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D4 = CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D5 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D6 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A1 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A2 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A4 = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A5 = CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A6 = 1'b1;
  assign RIOB33_X105Y143_IOB_X1Y143_O = CLBLM_L_X16Y136_SLICE_X23Y136_DQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A5 = 1'b1;
  assign RIOB33_X105Y143_IOB_X1Y144_O = CLBLM_R_X13Y138_SLICE_X19Y138_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_AX = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B1 = CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B2 = CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B3 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B4 = CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B5 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A6 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C2 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D6 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A1 = CLBLM_L_X16Y136_SLICE_X22Y136_AO5;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A2 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A3 = CLBLM_L_X16Y136_SLICE_X23Y136_AQ;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A4 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A5 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_A6 = CLBLM_R_X13Y136_SLICE_X19Y136_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B2 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B5 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_B6 = CLBLM_L_X16Y136_SLICE_X23Y136_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B4 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B5 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C1 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C2 = CLBLM_L_X16Y136_SLICE_X23Y136_CQ;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C4 = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C5 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_C6 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B6 = 1'b1;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_D = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_D = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D2 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D3 = CLBLM_L_X16Y136_SLICE_X23Y136_DQ;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D4 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D5 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_D6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y136_SLICE_X23Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A1 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A3 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A4 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A5 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_A6 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B1 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B2 = CLBLM_L_X16Y136_SLICE_X22Y136_BQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B3 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B5 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_B6 = CLBLM_L_X16Y136_SLICE_X22Y136_CO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C1 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C2 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C3 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C4 = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C5 = CLBLM_L_X16Y136_SLICE_X22Y136_DO6;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_C6 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D1 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D2 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D3 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D4 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D5 = 1'b1;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_D6 = CLBLM_R_X13Y137_SLICE_X19Y137_BQ;
  assign CLBLM_L_X16Y136_SLICE_X22Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A5 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A6 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A5 = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_AX = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B6 = CLBLM_R_X13Y149_SLICE_X18Y149_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign LIOB33_X0Y59_IOB_X0Y60_O = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign LIOB33_X0Y59_IOB_X0Y59_O = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C1 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A1 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A2 = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A4 = CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A5 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C1 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A6 = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C2 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_AX = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C3 = CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C2 = CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B1 = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B5 = CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B6 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C1 = CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C2 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C3 = CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C4 = CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C5 = CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C5 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C6 = 1'b1;
  assign RIOB33_X105Y145_IOB_X1Y145_O = CLBLM_L_X16Y138_SLICE_X22Y138_AQ;
  assign RIOB33_X105Y145_IOB_X1Y146_O = CLBLM_L_X16Y137_SLICE_X23Y137_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D1 = CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D2 = CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D3 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D4 = CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D5 = CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A2 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A3 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A4 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A5 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A6 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_AX = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A6 = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B2 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B3 = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B4 = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B5 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_BX = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C1 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C3 = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C4 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C5 = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D2 = CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_CX = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D1 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D2 = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D4 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D6 = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D4 = CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A2 = CLBLM_L_X16Y137_SLICE_X23Y137_BQ;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A3 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A4 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_A6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_DX = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D5 = CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D6 = CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B2 = CLBLM_L_X16Y137_SLICE_X23Y137_BQ;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B3 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B5 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_B6 = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C1 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C2 = CLBLM_L_X16Y137_SLICE_X23Y137_CQ;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C4 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C5 = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_C6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D1 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D2 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D3 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D4 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D5 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_D6 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X23Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A2 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A3 = CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A4 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A5 = CLBLM_L_X16Y137_SLICE_X23Y137_CQ;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_A6 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B3 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B4 = CLBLM_L_X16Y138_SLICE_X22Y138_AQ;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B5 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_B6 = 1'b1;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C1 = CLBLM_L_X16Y137_SLICE_X22Y137_AO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C2 = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C3 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C4 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_C6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D2 = CLBLM_L_X16Y137_SLICE_X23Y137_AO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D3 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D4 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D5 = CLBLM_L_X16Y137_SLICE_X22Y137_BO6;
  assign CLBLM_L_X16Y137_SLICE_X22Y137_D6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B1 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B2 = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign LIOB33_X0Y61_IOB_X0Y62_O = CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  assign LIOB33_X0Y61_IOB_X0Y61_O = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B3 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B6 = 1'b1;
  assign RIOB33_X105Y147_IOB_X1Y148_O = CLBLM_L_X16Y139_SLICE_X22Y139_BQ;
  assign RIOB33_X105Y147_IOB_X1Y147_O = CLBLM_L_X16Y137_SLICE_X23Y137_CQ;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A1 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A2 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_AX = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A5 = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A6 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B3 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B4 = CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B6 = CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C1 = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C2 = CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D2 = CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D3 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D4 = CLBLM_R_X5Y145_SLICE_X7Y145_AO5;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A2 = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A3 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A4 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A6 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_AX = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B2 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B4 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B5 = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B6 = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_BX = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C1 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C3 = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C4 = CLBLM_R_X3Y141_SLICE_X3Y141_CQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C6 = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CX = CLBLM_R_X3Y141_SLICE_X3Y141_CQ;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_A1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_A2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_A3 = CLBLM_L_X16Y138_SLICE_X23Y138_AQ;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_A4 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_A5 = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_A6 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D6 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_B1 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_B2 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_B3 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_B4 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_C1 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_B5 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_B6 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_C2 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_C3 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_C4 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_C5 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_C6 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_D1 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_D1 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_D2 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_D3 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_D4 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_D5 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_T1 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X23Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_A1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_A2 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_A3 = CLBLM_L_X16Y138_SLICE_X22Y138_AQ;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_A4 = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_A5 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_B1 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_B2 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_B3 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_B4 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_B5 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_B6 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_C1 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_C2 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_C3 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_C4 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_C5 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_C6 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_D1 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_D2 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_D3 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_D4 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_D5 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_D6 = 1'b1;
  assign CLBLM_L_X16Y138_SLICE_X22Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_D = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOB33_X0Y63_IOB_X0Y63_O = 1'b1;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_D = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A6 = LIOB33_X0Y189_IOB_X0Y190_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_AX = LIOB33_X0Y193_IOB_X0Y194_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B6 = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A1 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A2 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_BX = LIOB33_X0Y195_IOB_X0Y195_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A3 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C6 = LIOB33_X0Y191_IOB_X0Y192_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_CE = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B1 = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B3 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_CX = LIOB33_X0Y195_IOB_X0Y196_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B6 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D6 = LIOB33_X0Y193_IOB_X0Y193_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C4 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_DX = LIOB33_X0Y197_IOB_X0Y197_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D2 = CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D6 = CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_AX = 1'b0;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A1 = CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A2 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A3 = CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A4 = CLBLL_L_X2Y153_SLICE_X0Y153_BQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A5 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_AX = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B1 = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B2 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B3 = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B4 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B5 = CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B6 = CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_BX = 1'b0;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_BX = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C1 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C3 = CLBLL_L_X2Y153_SLICE_X1Y153_BQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C4 = CLBLL_L_X2Y153_SLICE_X0Y153_CQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C5 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C6 = CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_CE = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_CIN = CLBLM_R_X5Y143_SLICE_X6Y143_COUT;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_CX = 1'b0;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D3 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_A1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D1 = CLBLL_L_X2Y152_SLICE_X0Y152_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D6 = CLBLL_L_X2Y153_SLICE_X0Y153_BQ;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_A2 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_A3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_A4 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_A5 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_B5 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_B6 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_B1 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_B2 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_B3 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_B4 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_C3 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_C4 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_C5 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_C6 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_C1 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_C2 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_D1 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_D2 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_D3 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_D4 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_D5 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X23Y139_D6 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_A1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_A2 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_A3 = CLBLM_L_X16Y139_SLICE_X22Y139_AQ;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_A4 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_A5 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_A6 = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_B2 = CLBLM_L_X16Y139_SLICE_X22Y139_BQ;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_B3 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_B5 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_B6 = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_C1 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_C2 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_C3 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_C4 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_C5 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_C6 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_D1 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_D2 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_D3 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_D4 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_D5 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_D6 = 1'b1;
  assign CLBLM_L_X16Y139_SLICE_X22Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLL_L_X4Y135_SLICE_X4Y135_B5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A1 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A2 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A3 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A4 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A6 = 1'b1;
  assign RIOB33_X105Y139_IOB_X1Y140_O = CLBLM_L_X16Y139_SLICE_X22Y139_AQ;
  assign RIOB33_X105Y139_IOB_X1Y139_O = CLBLM_L_X16Y138_SLICE_X23Y138_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A6 = 1'b1;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_D = LIOB33_X0Y195_IOB_X0Y196_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B1 = CLBLM_R_X13Y129_SLICE_X18Y129_B5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B2 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B3 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_D = LIOB33_X0Y195_IOB_X0Y195_I;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B4 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B5 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_A1 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_A2 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_A3 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_A4 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_A5 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_A6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_B6 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_B1 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_B2 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_B3 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_B4 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_B5 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_B6 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_C1 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_C2 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_C3 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_C4 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_C5 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_C6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C1 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C2 = CLBLM_R_X13Y129_SLICE_X18Y129_CQ;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_D1 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_D2 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_D3 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_D4 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_D5 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X23Y140_D6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C3 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_DQ;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_A1 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_A2 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_A3 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_A4 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_A5 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_A6 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_AX = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_CE = CLBLM_R_X13Y129_SLICE_X19Y129_CO6;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_B1 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_B2 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_B3 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_B4 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_B5 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_B6 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_BX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_C1 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_C2 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_C3 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_C4 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_C5 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_C6 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_CE = CLBLM_L_X16Y143_SLICE_X22Y143_AO6;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_B4 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_CX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_B5 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_D1 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_D2 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_D3 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_D4 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_D5 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_D6 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_B6 = CLBLM_R_X15Y148_SLICE_X21Y148_CO6;
  assign LIOI3_X0Y53_OLOGIC_X0Y54_T1 = 1'b1;
  assign CLBLM_L_X16Y140_SLICE_X22Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y58_T1 = 1'b1;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_B5Q;
  assign LIOI3_X0Y53_OLOGIC_X0Y53_T1 = 1'b1;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_C3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D5 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_C4 = CLBLM_R_X15Y148_SLICE_X21Y148_AO5;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_C5 = CLBLM_R_X15Y148_SLICE_X21Y148_DO6;
  assign CLBLM_R_X15Y148_SLICE_X21Y148_C6 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A1 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A3 = CLBLL_L_X2Y158_SLICE_X1Y158_AQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A4 = CLBLL_L_X2Y156_SLICE_X0Y156_AO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A5 = CLBLL_L_X2Y158_SLICE_X1Y158_DQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A6 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_AX = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B1 = CLBLL_L_X2Y156_SLICE_X0Y156_DO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B2 = CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B3 = CLBLL_L_X2Y155_SLICE_X0Y155_AQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B4 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B5 = CLBLL_L_X2Y158_SLICE_X1Y158_AQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B6 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_BX = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C1 = CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C2 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C3 = CLBLL_L_X2Y158_SLICE_X1Y158_BQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C4 = CLBLL_L_X2Y155_SLICE_X0Y155_BQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C5 = CLBLL_L_X2Y157_SLICE_X0Y157_DO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C6 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A6 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C6 = 1'b1;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_D = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D6 = 1'b1;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_D = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A2 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A3 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_AX = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B1 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C6 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C1 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C2 = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_A1 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_A2 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_A3 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_A4 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_A5 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_A6 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_AX = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_B1 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_B2 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_B3 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_B4 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_B5 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_B6 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_BX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_C1 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_C2 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_C3 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_C4 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_C5 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_C6 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_CE = CLBLM_L_X16Y142_SLICE_X22Y142_CO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B6 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_CX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_D1 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_D2 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_D3 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_D4 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_D5 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_D6 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_DX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_L_X16Y141_SLICE_X23Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_A1 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_A2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_A3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_A5 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_A6 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_AX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_B2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_B3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_B4 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_B5 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_B6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_BX = CLBLM_R_X15Y140_SLICE_X21Y140_AO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_C1 = CLBLM_R_X15Y141_SLICE_X20Y141_CQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_C2 = CLBLM_L_X16Y141_SLICE_X22Y141_AQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_C3 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_C5 = CLBLM_R_X15Y141_SLICE_X21Y141_CQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_C6 = CLBLM_L_X16Y141_SLICE_X23Y141_BQ;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_CE = CLBLM_L_X16Y141_SLICE_X22Y141_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D4 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D5 = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_CX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_D1 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_D2 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_D3 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_D4 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_D5 = 1'b1;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_D6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D6 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X16Y141_SLICE_X22Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A1 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A2 = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A4 = CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A3 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A5 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A6 = CLBLM_R_X13Y150_SLICE_X18Y150_CO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B6 = CLBLM_R_X13Y144_SLICE_X19Y144_CO5;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_A1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_A2 = CLBLL_L_X2Y156_SLICE_X0Y156_BQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_A3 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_A4 = CLBLL_L_X2Y156_SLICE_X0Y156_CQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_A5 = CLBLL_L_X2Y155_SLICE_X0Y155_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_A6 = CLBLL_L_X2Y156_SLICE_X0Y156_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_AX = CLBLL_L_X2Y158_SLICE_X1Y158_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_B2 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_B3 = CLBLL_L_X2Y158_SLICE_X1Y158_DQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_B4 = CLBLL_L_X2Y158_SLICE_X0Y158_BQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_B5 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_B6 = CLBLL_L_X2Y156_SLICE_X0Y156_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_BX = CLBLL_L_X2Y158_SLICE_X1Y158_DQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_C1 = CLBLL_L_X2Y158_SLICE_X1Y158_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_C2 = CLBLL_L_X2Y155_SLICE_X0Y155_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_C3 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_C4 = CLBLL_L_X2Y156_SLICE_X0Y156_BQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_C5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_C6 = CLBLL_L_X2Y156_SLICE_X0Y156_CQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A1 = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A2 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A3 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A5 = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_CX = CLBLL_L_X2Y158_SLICE_X0Y158_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A6 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_D1 = CLBLL_L_X2Y156_SLICE_X0Y156_BQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_D2 = CLBLL_L_X2Y156_SLICE_X0Y156_CQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_D3 = CLBLL_L_X2Y156_SLICE_X0Y156_DQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_D4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_D6 = CLBLL_L_X2Y156_SLICE_X0Y156_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_DX = CLBLL_L_X2Y155_SLICE_X0Y155_AQ;
  assign CLBLL_L_X2Y156_SLICE_X0Y156_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B2 = CLBLM_R_X5Y147_SLICE_X6Y147_BO5;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B3 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_A1 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_A2 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_A3 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_A4 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_A5 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_A6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A1 = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A2 = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_B1 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_B2 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_B3 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_B4 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_B5 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_B6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A6 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_C1 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_C2 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_C3 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_C4 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_C5 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_C6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C1 = CLBLM_R_X5Y151_SLICE_X7Y151_AO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C2 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C3 = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_D1 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_D2 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_D3 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_D4 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_D5 = 1'b1;
  assign CLBLL_L_X2Y156_SLICE_X1Y156_D6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D2 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D3 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_A1 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_A2 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_A3 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_A4 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_A5 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_A6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D6 = CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_AX = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_B1 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_B2 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_B3 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_B4 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_B5 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_B6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D6 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_C1 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_C2 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_C3 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_C4 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_C5 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_C6 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_CE = CLBLM_L_X16Y141_SLICE_X22Y141_AO6;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_D1 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_D2 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_D3 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_D4 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_D5 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_D6 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X23Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_A1 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_A4 = CLBLM_R_X15Y142_SLICE_X21Y142_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_A5 = CLBLM_L_X16Y142_SLICE_X23Y142_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_A6 = 1'b1;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_AX = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_B1 = CLBLM_R_X15Y144_SLICE_X21Y144_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_B2 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_B3 = CLBLM_L_X16Y142_SLICE_X22Y142_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_B4 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_B5 = CLBLM_L_X16Y142_SLICE_X22Y142_AO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_BX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_C1 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_C2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_C3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_C5 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_C6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_CE = CLBLM_L_X16Y142_SLICE_X22Y142_CO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_CX = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_D1 = CLBLM_L_X16Y142_SLICE_X23Y142_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_D3 = CLBLM_L_X16Y142_SLICE_X22Y142_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_D4 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_D5 = CLBLM_R_X15Y144_SLICE_X21Y144_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_D6 = CLBLM_R_X15Y142_SLICE_X21Y142_AQ;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_DX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_L_X16Y142_SLICE_X22Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A6 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A1 = CLBLL_L_X2Y157_SLICE_X0Y157_BO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A3 = CLBLL_L_X2Y158_SLICE_X1Y158_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A4 = CLBLL_L_X2Y158_SLICE_X0Y158_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A5 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_A6 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_D1 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_AX = CLBLL_L_X2Y158_SLICE_X1Y158_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B1 = CLBLL_L_X2Y155_SLICE_X0Y155_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B2 = CLBLL_L_X2Y157_SLICE_X0Y157_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B3 = CLBLL_L_X2Y157_SLICE_X0Y157_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B4 = CLBLL_L_X2Y157_SLICE_X0Y157_CQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_B6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign LIOI3_X0Y55_OLOGIC_X0Y56_T1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_BX = CLBLL_L_X2Y158_SLICE_X0Y158_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C2 = CLBLL_L_X2Y157_SLICE_X0Y157_CQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C3 = CLBLL_L_X2Y155_SLICE_X0Y155_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C5 = CLBLL_L_X2Y157_SLICE_X0Y157_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_C6 = CLBLL_L_X2Y158_SLICE_X1Y158_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_D1 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A1 = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A2 = CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_CX = CLBLL_L_X2Y158_SLICE_X0Y158_DQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D2 = CLBLL_L_X2Y157_SLICE_X0Y157_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D3 = CLBLL_L_X2Y157_SLICE_X0Y157_DQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D4 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D5 = CLBLL_L_X2Y157_SLICE_X0Y157_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_D6 = CLBLL_L_X2Y157_SLICE_X0Y157_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A6 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_DX = CLBLL_L_X2Y155_SLICE_X0Y155_BQ;
  assign CLBLL_L_X2Y157_SLICE_X0Y157_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B3 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B5 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C1 = CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C3 = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C4 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C5 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C6 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D2 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D3 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_A6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D6 = CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A1 = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_B6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A6 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_C6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B1 = CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B2 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B3 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B4 = CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B5 = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B6 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D1 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D2 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D3 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D4 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D5 = 1'b1;
  assign CLBLL_L_X2Y157_SLICE_X1Y157_D6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C6 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D2 = CLBLM_R_X5Y148_SLICE_X7Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D3 = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D4 = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D5 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D6 = CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_A1 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_A2 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_A3 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_A4 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_A5 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_A6 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_B1 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_B2 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_B3 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_B4 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_B5 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_B6 = 1'b1;
  assign LIOI3_X0Y51_OLOGIC_X0Y52_T1 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_C1 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_C2 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_C3 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_C4 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_C5 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_C6 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_D1 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_D2 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_D3 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_D4 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_D5 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X23Y143_D6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D3 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_A1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_A3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_A4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_A5 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_D = LIOB33_X0Y177_IOB_X0Y178_I;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_AX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B5 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_B1 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_B2 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_B3 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_B4 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_B5 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_B6 = 1'b1;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_D = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_BX = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_C1 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_C2 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_C3 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_C4 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_C5 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_C6 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_CE = CLBLM_L_X16Y143_SLICE_X22Y143_AO6;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_CX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_D1 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_D2 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_D3 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_D4 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_D5 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_D6 = 1'b1;
  assign CLBLM_L_X16Y143_SLICE_X22Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y51_OLOGIC_X0Y51_T1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D4 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_A6 = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_AX = LIOB33_X0Y179_IOB_X0Y180_I;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B1 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B2 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B3 = CLBLL_L_X2Y158_SLICE_X0Y158_AQ;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B4 = CLBLL_L_X2Y158_SLICE_X0Y158_DQ;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_B6 = CLBLL_L_X2Y157_SLICE_X0Y157_CO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_BX = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_C6 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_CX = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_D6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A1 = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A2 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_DX = LIOB33_X0Y177_IOB_X0Y178_I;
  assign CLBLL_L_X2Y158_SLICE_X0Y158_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A3 = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A4 = CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A5 = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A6 = CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C5 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C6 = CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_A6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D1 = CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_AX = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_B6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_BX = LIOB33_X0Y161_IOB_X0Y162_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_C6 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_CE = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A6 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B1 = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B2 = CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B3 = CLBLM_L_X16Y142_SLICE_X22Y142_AO5;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_CX = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B4 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D1 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D2 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D3 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D4 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D5 = 1'b1;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_D6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_DX = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLL_L_X2Y158_SLICE_X1Y158_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C5 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D3 = CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D6 = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C4 = CLBLL_L_X26Y133_SLICE_X38Y133_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C6 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOB33_X105Y141_IOB_X1Y142_O = CLBLM_R_X13Y138_SLICE_X19Y138_BQ;
  assign RIOB33_X105Y141_IOB_X1Y141_O = CLBLM_R_X13Y138_SLICE_X19Y138_AQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B3 = CLBLM_R_X15Y128_SLICE_X20Y128_CQ;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_B4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A1 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A2 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A3 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A5 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_A6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B1 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B2 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B3 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B5 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_B6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C1 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C2 = CLBLM_R_X15Y128_SLICE_X20Y128_CQ;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C1 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C2 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C3 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C5 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_C6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C3 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D1 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D2 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D3 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D5 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X19Y128_D6 = 1'b1;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_C6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A1 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A2 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A3 = CLBLM_R_X13Y128_SLICE_X18Y128_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A4 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A5 = CLBLM_R_X13Y128_SLICE_X18Y128_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A1 = CLBLM_R_X5Y150_SLICE_X7Y150_DO5;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A2 = CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A3 = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A4 = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A5 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A6 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B1 = CLBLM_R_X13Y128_SLICE_X18Y128_B5Q;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B2 = CLBLM_R_X13Y128_SLICE_X18Y128_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B4 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B5 = CLBLM_R_X13Y128_SLICE_X18Y128_A5Q;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_B6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C1 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C5 = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_C5 = CLBLM_R_X13Y128_SLICE_X18Y128_B5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_CE = CLBLM_L_X12Y129_SLICE_X17Y129_CO6;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D1 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D6 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D3 = 1'b1;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_D4 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y128_SLICE_X18Y128_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y128_SLICE_X20Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A3 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B1 = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B3 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B4 = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B6 = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C1 = CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C2 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C5 = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C6 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D4 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D5 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D6 = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_D1 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign LIOI3_X0Y59_OLOGIC_X0Y60_T1 = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_D1 = CLBLM_L_X12Y128_SLICE_X16Y128_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C4 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_T1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C5 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B3 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A2 = CLBLM_R_X13Y130_SLICE_X18Y130_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A3 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A4 = CLBLM_R_X13Y129_SLICE_X19Y129_BO6;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A5 = CLBLM_R_X15Y129_SLICE_X20Y129_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B4 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_A6 = 1'b1;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_D = LIOB33_X0Y179_IOB_X0Y180_I;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B1 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B3 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B4 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B5 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_B6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C1 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C3 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C4 = CLBLM_R_X13Y136_SLICE_X19Y136_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C5 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_C6 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D1 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_BX = 1'b0;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D3 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D4 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D5 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_D6 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X19Y129_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C1 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A1 = CLBLM_R_X13Y129_SLICE_X18Y129_B5Q;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A2 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C2 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A3 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A4 = CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_A5 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D3 = CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A3 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A5 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C3 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D5 = CLBLM_L_X16Y136_SLICE_X22Y136_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B3 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B4 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D6 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C6 = CLBLM_L_X12Y132_SLICE_X17Y132_A5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C1 = CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C2 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C5 = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C6 = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C4 = 1'b1;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C5 = CLBLM_R_X13Y129_SLICE_X18Y129_B5Q;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_C6 = CLBLM_R_X13Y129_SLICE_X18Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D1 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D2 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D6 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D3 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D4 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_D6 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y129_SLICE_X18Y129_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C5 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D3 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D6 = CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D6 = CLBLM_L_X12Y131_SLICE_X17Y131_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B1 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B2 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B3 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B2 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B6 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D5 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D6 = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A1 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A2 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A3 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A4 = CLBLM_R_X13Y130_SLICE_X19Y130_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A5 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_A6 = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B1 = CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B2 = CLBLM_L_X16Y136_SLICE_X22Y136_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B3 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B4 = CLBLM_R_X13Y136_SLICE_X19Y136_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B5 = CLBLM_R_X15Y130_SLICE_X20Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_B6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C1 = CLBLM_L_X16Y136_SLICE_X22Y136_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C2 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C3 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C5 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_C6 = CLBLM_R_X13Y136_SLICE_X19Y136_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B1 = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B2 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B3 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D2 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D3 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D4 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D5 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_D6 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X19Y130_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A1 = CLBLM_R_X13Y129_SLICE_X19Y129_BO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A2 = 1'b1;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A3 = CLBLM_L_X12Y129_SLICE_X17Y129_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A4 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_A6 = CLBLM_L_X12Y130_SLICE_X17Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B1 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B2 = CLBLM_R_X13Y136_SLICE_X19Y136_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B3 = CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B4 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B5 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_B6 = CLBLM_R_X13Y129_SLICE_X18Y129_CQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C1 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C3 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C4 = CLBLM_R_X13Y129_SLICE_X18Y129_CQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C5 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_C6 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_CE = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D1 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D2 = CLBLM_R_X13Y130_SLICE_X19Y130_CO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D3 = CLBLM_R_X13Y129_SLICE_X19Y129_BO5;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D4 = CLBLM_R_X13Y129_SLICE_X18Y129_CQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D5 = CLBLM_R_X13Y129_SLICE_X18Y129_BQ;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_D6 = CLBLM_R_X13Y129_SLICE_X19Y129_DO6;
  assign CLBLM_R_X13Y130_SLICE_X18Y130_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_D1 = CLBLL_L_X2Y116_SLICE_X0Y116_AQ;
  assign LIOI3_X0Y61_OLOGIC_X0Y62_T1 = 1'b1;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_D1 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign LIOI3_X0Y61_OLOGIC_X0Y61_T1 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A1 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A2 = CLBLM_R_X13Y130_SLICE_X18Y130_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A3 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A4 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A5 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_A6 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B1 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B2 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B3 = CLBLM_R_X13Y131_SLICE_X19Y131_CQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B4 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B5 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_B6 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C1 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C2 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C3 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C4 = CLBLM_R_X13Y131_SLICE_X19Y131_DQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C5 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_C6 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_CE = CLBLM_R_X13Y130_SLICE_X18Y130_DO6;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D1 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D2 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D3 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D4 = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D5 = CLBLM_R_X13Y132_SLICE_X18Y132_DQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_D6 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X13Y131_SLICE_X19Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A1 = CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A2 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A3 = CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A4 = CLBLM_R_X13Y131_SLICE_X18Y131_BO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A5 = CLBLM_R_X13Y131_SLICE_X18Y131_CO6;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_A6 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_AX = CLBLM_R_X15Y131_SLICE_X20Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B1 = CLBLM_L_X12Y131_SLICE_X16Y131_A5Q;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B2 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B3 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B4 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B5 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_B6 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_BX = CLBLM_R_X13Y131_SLICE_X19Y131_BQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C2 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C4 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C5 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_C6 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_CE = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_CX = CLBLM_R_X13Y131_SLICE_X19Y131_DQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D1 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D2 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D3 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D4 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D5 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_D6 = 1'b1;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_DX = CLBLM_R_X13Y131_SLICE_X19Y131_AQ;
  assign CLBLM_R_X13Y131_SLICE_X18Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_D = LIOB33_X0Y183_IOB_X0Y184_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_D = LIOB33_X0Y183_IOB_X0Y183_I;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = CLBLM_L_X16Y139_SLICE_X22Y139_AQ;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_B6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_C6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D2 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D3 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X19Y132_D6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A2 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A3 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A4 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A5 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B1 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B2 = CLBLM_R_X13Y138_SLICE_X18Y138_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B3 = CLBLM_L_X12Y131_SLICE_X17Y131_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B5 = CLBLM_R_X13Y134_SLICE_X19Y134_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_B6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C1 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C4 = CLBLM_L_X12Y131_SLICE_X17Y131_A5Q;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C5 = CLBLM_L_X12Y132_SLICE_X17Y132_A5Q;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_C6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D1 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D2 = CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D3 = CLBLM_R_X13Y135_SLICE_X19Y135_DQ;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D4 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D5 = CLBLM_R_X13Y132_SLICE_X18Y132_D5Q;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_D6 = 1'b1;
  assign CLBLM_R_X13Y132_SLICE_X18Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B3 = CLBLM_R_X15Y129_SLICE_X20Y129_CQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_B4 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A1 = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A2 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A3 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A4 = CLBLM_R_X15Y134_SLICE_X21Y134_BQ;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A5 = CLBLM_R_X15Y133_SLICE_X21Y133_AQ;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B2 = CLBLM_R_X15Y133_SLICE_X21Y133_BQ;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B3 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B4 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B5 = CLBLM_R_X15Y133_SLICE_X21Y133_CQ;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C3 = CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C5 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_CE = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C1 = CLBLM_R_X15Y131_SLICE_X20Y131_AQ;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C2 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_C3 = CLBLM_R_X13Y130_SLICE_X19Y130_AQ;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D1 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D2 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D3 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D4 = CLBLM_R_X13Y136_SLICE_X19Y136_AQ;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D6 = CLBLM_L_X16Y136_SLICE_X23Y136_AQ;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A1 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A3 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A4 = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A5 = CLBLM_R_X13Y133_SLICE_X19Y133_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B1 = CLBLM_R_X13Y136_SLICE_X18Y136_B5Q;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B2 = CLBLM_R_X13Y133_SLICE_X19Y133_B5Q;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B4 = CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B5 = CLBLM_L_X12Y138_SLICE_X17Y138_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C1 = CLBLM_R_X15Y134_SLICE_X21Y134_BQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C2 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C3 = CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C4 = CLBLM_R_X13Y132_SLICE_X18Y132_CO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C6 = CLBLM_R_X15Y136_SLICE_X21Y136_CQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D3 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = CLBLM_L_X16Y136_SLICE_X23Y136_CQ;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_A5Q;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D4 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = CLBLM_L_X16Y136_SLICE_X23Y136_BQ;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_A1 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_A2 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_A3 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_A4 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_A5 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_A6 = 1'b1;
  assign CLBLM_R_X15Y129_SLICE_X20Y129_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_B1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_B2 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_B3 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_B4 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_B5 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_B6 = 1'b1;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_C1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_C3 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_C4 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_C5 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_C6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_D1 = CLBLM_R_X15Y152_SLICE_X21Y152_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_D2 = 1'b1;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_D3 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_D4 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_D5 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y150_SLICE_X23Y150_D6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A2 = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A3 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A4 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A5 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A6 = 1'b1;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_A2 = 1'b1;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_A3 = CLBLM_R_X15Y152_SLICE_X21Y152_AQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_A4 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_A6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B1 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B2 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_AX = 1'b0;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B3 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_B2 = CLBLM_L_X16Y150_SLICE_X23Y150_DO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_B3 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_B4 = CLBLM_R_X15Y151_SLICE_X21Y151_A5Q;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_B6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C1 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C2 = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_BX = CLBLM_L_X16Y150_SLICE_X23Y150_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_C1 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_C2 = CLBLM_L_X16Y150_SLICE_X23Y150_AO5;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_C3 = CLBLM_R_X15Y150_SLICE_X21Y150_DO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_C4 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_C6 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D6 = 1'b1;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_CX = CLBLM_R_X15Y150_SLICE_X21Y150_DO6;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_D = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_D1 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_D2 = CLBLM_L_X16Y150_SLICE_X23Y150_CO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_D3 = CLBLM_L_X16Y150_SLICE_X23Y150_BO5;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_D4 = CLBLM_R_X15Y152_SLICE_X21Y152_BQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_D5 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_D6 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A2 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_DX = CLBLM_L_X16Y150_SLICE_X23Y150_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A4 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A5 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B1 = CLBLM_L_X12Y130_SLICE_X16Y130_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B2 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B4 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B5 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B6 = CLBLM_L_X12Y130_SLICE_X17Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C5 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A1 = CLBLM_R_X15Y135_SLICE_X21Y135_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A2 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A3 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A5 = CLBLM_R_X15Y134_SLICE_X21Y134_AQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B1 = CLBLM_R_X15Y134_SLICE_X21Y134_CQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B2 = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B3 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B4 = CLBLM_R_X15Y135_SLICE_X21Y135_AQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B5 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B4 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C1 = CLBLM_R_X15Y133_SLICE_X21Y133_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C2 = CLBLM_R_X13Y135_SLICE_X19Y135_CQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C3 = CLBLM_R_X13Y132_SLICE_X18Y132_BO5;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C4 = CLBLM_R_X15Y136_SLICE_X21Y136_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C6 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_CE = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D1 = CLBLM_R_X15Y133_SLICE_X21Y133_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D2 = CLBLM_R_X15Y136_SLICE_X21Y136_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D3 = CLBLM_R_X15Y135_SLICE_X21Y135_CO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D4 = CLBLM_R_X15Y135_SLICE_X21Y135_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D5 = CLBLM_R_X13Y135_SLICE_X19Y135_DO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D6 = CLBLM_R_X15Y133_SLICE_X21Y133_CQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A1 = CLBLM_R_X13Y133_SLICE_X19Y133_A5Q;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A2 = CLBLM_R_X13Y136_SLICE_X18Y136_A5Q;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A4 = CLBLM_R_X13Y136_SLICE_X18Y136_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A5 = CLBLM_R_X13Y133_SLICE_X19Y133_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C1 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B1 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B2 = CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C2 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B3 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B4 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B5 = CLBLM_R_X15Y137_SLICE_X20Y137_D_CY;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D3 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C4 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C1 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C2 = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C3 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C4 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C5 = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C6 = CLBLM_L_X12Y131_SLICE_X16Y131_A5Q;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D1 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D2 = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D3 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D4 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D5 = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_A6 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D3 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A2 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A4 = CLBLM_R_X15Y152_SLICE_X21Y152_BQ;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A5 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_A6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_AX = CLBLM_L_X16Y152_SLICE_X23Y152_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B3 = CLBLM_L_X16Y151_SLICE_X23Y151_AQ;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B4 = CLBLM_L_X16Y150_SLICE_X23Y150_BO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_B6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D6 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C1 = CLBLM_L_X16Y150_SLICE_X23Y150_AO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C2 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C3 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C4 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C5 = CLBLM_R_X15Y152_SLICE_X20Y152_AQ;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_C6 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_B4 = CLBLM_R_X15Y152_SLICE_X20Y152_BO6;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D2 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D3 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D4 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D5 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_D6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A1 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A2 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X16Y151_SLICE_X23Y151_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A3 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A4 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A5 = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A1 = CLBLM_R_X15Y152_SLICE_X20Y152_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A2 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A3 = CLBLM_L_X16Y151_SLICE_X23Y151_AO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A4 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A5 = CLBLM_L_X16Y150_SLICE_X23Y150_AO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_A6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A6 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B1 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_AX = CLBLM_L_X16Y151_SLICE_X23Y151_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B1 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B2 = CLBLM_L_X16Y150_SLICE_X23Y150_BO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B3 = CLBLM_L_X16Y151_SLICE_X23Y151_CO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B4 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B5 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_B6 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C1 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_BX = CLBLM_L_X16Y151_SLICE_X23Y151_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C1 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C2 = CLBLM_L_X16Y151_SLICE_X23Y151_BO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C3 = CLBLM_R_X15Y151_SLICE_X20Y151_BQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C4 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C5 = CLBLM_R_X15Y151_SLICE_X21Y151_CO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_C6 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_CIN = CLBLM_L_X16Y150_SLICE_X22Y150_COUT;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D2 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D3 = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D4 = CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D5 = CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_CX = CLBLM_L_X16Y151_SLICE_X23Y151_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D6 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D1 = 1'b1;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D2 = CLBLM_R_X15Y151_SLICE_X20Y151_BQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D3 = CLBLM_R_X15Y151_SLICE_X21Y151_CO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D4 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_D6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A1 = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X16Y151_SLICE_X22Y151_DX = 1'b0;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A2 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A3 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A4 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A5 = CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A6 = CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B1 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B2 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B4 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B5 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B6 = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C2 = CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C3 = CLBLM_L_X12Y132_SLICE_X17Y132_B5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C5 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C6 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D2 = CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D3 = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D6 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B2 = CLBLM_R_X13Y146_SLICE_X19Y146_AO5;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A1 = CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A2 = CLBLM_R_X15Y136_SLICE_X21Y136_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A3 = CLBLM_R_X13Y135_SLICE_X19Y135_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A4 = CLBLM_R_X15Y133_SLICE_X21Y133_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A5 = CLBLM_R_X13Y132_SLICE_X18Y132_AO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_D5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_AX = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B1 = CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B2 = CLBLM_R_X13Y135_SLICE_X19Y135_BQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B4 = CLBLM_R_X15Y134_SLICE_X21Y134_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B5 = CLBLM_R_X15Y137_SLICE_X21Y137_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B6 = CLBLM_R_X13Y133_SLICE_X18Y133_AO5;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_D6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_BX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C2 = CLBLM_R_X13Y136_SLICE_X19Y136_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C3 = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C4 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C5 = CLBLM_R_X15Y134_SLICE_X20Y134_DQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C6 = CLBLL_L_X26Y135_SLICE_X38Y135_AO5;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_CE = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_CX = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D1 = CLBLM_R_X15Y133_SLICE_X21Y133_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D2 = CLBLM_R_X15Y134_SLICE_X21Y134_CQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D3 = CLBLM_R_X15Y137_SLICE_X21Y137_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D5 = CLBLM_R_X15Y138_SLICE_X21Y138_AQ;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D6 = 1'b1;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_DX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A1 = CLBLM_R_X13Y138_SLICE_X18Y138_A5Q;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A2 = CLBLM_R_X13Y134_SLICE_X19Y134_A5Q;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A4 = CLBLM_L_X12Y138_SLICE_X17Y138_BQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A5 = CLBLM_R_X13Y134_SLICE_X19Y134_B5Q;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_AX = CLBLM_R_X15Y143_SLICE_X21Y143_AO5;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B2 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B3 = CLBLM_R_X13Y135_SLICE_X19Y135_AO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B4 = CLBLM_L_X16Y135_SLICE_X22Y135_CO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B5 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B6 = CLBLM_R_X13Y135_SLICE_X18Y135_CO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_BX = CLBLM_L_X16Y136_SLICE_X22Y136_AO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C1 = CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C2 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C3 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C4 = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C5 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C6 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_CE = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D1 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D4 = CLBLM_R_X15Y135_SLICE_X21Y135_BQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D5 = CLBLM_R_X13Y135_SLICE_X19Y135_DQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D6 = CLBLM_R_X15Y138_SLICE_X21Y138_BQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B3 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A1 = CLBLM_L_X16Y152_SLICE_X22Y152_A_XOR;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A2 = CLBLM_R_X15Y152_SLICE_X20Y152_DO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A3 = CLBLM_L_X16Y152_SLICE_X23Y152_AQ;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A4 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A5 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_A6 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B1 = CLBLM_L_X16Y154_SLICE_X22Y154_A_CY;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B2 = CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B3 = CLBLM_L_X16Y153_SLICE_X22Y153_C_XOR;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B4 = CLBLM_L_X16Y153_SLICE_X23Y153_BO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B5 = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_B6 = CLBLM_L_X16Y153_SLICE_X23Y153_AO5;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C1 = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C2 = CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C3 = CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C4 = CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_C6 = CLBLM_L_X16Y153_SLICE_X23Y153_BO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D1 = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D2 = CLBLM_R_X15Y152_SLICE_X21Y152_DO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D3 = CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D4 = CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_D6 = CLBLM_L_X16Y150_SLICE_X22Y150_A_XOR;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = CLBLM_R_X11Y133_SLICE_X15Y133_A_CY;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = CLBLM_R_X11Y133_SLICE_X14Y133_D_CY;
  assign CLBLM_L_X16Y152_SLICE_X23Y152_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A1 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A2 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A4 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A5 = CLBLM_L_X16Y152_SLICE_X23Y152_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_A6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B1 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B2 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B3 = CLBLM_L_X16Y150_SLICE_X22Y150_A_XOR;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B4 = CLBLM_R_X15Y152_SLICE_X21Y152_DO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_B6 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = CLBLM_L_X12Y131_SLICE_X16Y131_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_BX = CLBLM_L_X16Y152_SLICE_X23Y152_DO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C4 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C5 = CLBLM_L_X16Y150_SLICE_X23Y150_AO5;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_C6 = CLBLM_R_X15Y151_SLICE_X21Y151_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = CLBLM_L_X12Y132_SLICE_X17Y132_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_CX = CLBLM_R_X15Y152_SLICE_X21Y152_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X2Y139_SLICE_X1Y139_DO5;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D1 = CLBLM_R_X15Y150_SLICE_X21Y150_CO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D2 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D3 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D4 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D5 = 1'b1;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_D6 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_DX = CLBLM_R_X15Y150_SLICE_X21Y150_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = CLBLM_L_X12Y131_SLICE_X16Y131_A5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = CLBLM_R_X15Y128_SLICE_X20Y128_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A1 = CLBLM_R_X13Y136_SLICE_X19Y136_AQ;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A3 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A4 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A5 = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A6 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B5 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B1 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B2 = CLBLM_R_X13Y136_SLICE_X19Y136_BQ;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B5 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B6 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C1 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C2 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C3 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C4 = CLBLM_R_X13Y136_SLICE_X19Y136_BQ;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C5 = CLBLM_R_X13Y137_SLICE_X19Y137_BQ;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C6 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_D = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_D = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D1 = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D2 = CLBLM_R_X15Y131_SLICE_X21Y131_BO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D3 = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D4 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D5 = CLBLM_L_X12Y129_SLICE_X16Y129_BQ;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D6 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A1 = CLBLM_R_X15Y136_SLICE_X21Y136_CQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A2 = CLBLM_R_X15Y136_SLICE_X21Y136_AQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A3 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A5 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B1 = CLBLM_R_X15Y136_SLICE_X21Y136_DQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B2 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B3 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B4 = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B5 = CLBLM_R_X15Y136_SLICE_X21Y136_BQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C1 = CLBLM_R_X15Y136_SLICE_X21Y136_DQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C2 = CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C4 = CLBLM_R_X15Y133_SLICE_X21Y133_CQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C5 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C6 = CLBLM_R_X13Y132_SLICE_X18Y132_CO5;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_CE = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D2 = CLBLM_R_X13Y138_SLICE_X18Y138_CO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D3 = CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D4 = CLBLM_R_X13Y136_SLICE_X18Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D6 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A1 = CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A2 = CLBLM_L_X16Y151_SLICE_X22Y151_D_XOR;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A3 = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_A6 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B3 = CLBLM_L_X16Y151_SLICE_X23Y151_AQ;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B4 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B5 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_B6 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_C6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B6 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X23Y153_D6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A1 = CLBLM_L_X12Y132_SLICE_X17Y132_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A2 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A4 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A5 = CLBLM_L_X12Y132_SLICE_X17Y132_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A6 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A1 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A2 = CLBLM_R_X15Y152_SLICE_X21Y152_BQ;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A3 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A4 = CLBLM_L_X16Y150_SLICE_X22Y150_D_XOR;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A5 = CLBLM_L_X16Y150_SLICE_X23Y150_AO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_A6 = CLBLM_R_X15Y153_SLICE_X21Y153_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_AX = CLBLM_R_X15Y153_SLICE_X21Y153_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B1 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B2 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B3 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B4 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B5 = CLBLM_R_X15Y152_SLICE_X20Y152_AO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_B6 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_BX = CLBLM_R_X15Y152_SLICE_X20Y152_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C3 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C1 = CLBLM_L_X16Y151_SLICE_X23Y151_AQ;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C2 = CLBLM_L_X16Y153_SLICE_X23Y153_AO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C3 = CLBLM_L_X16Y151_SLICE_X22Y151_B_XOR;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C4 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C5 = CLBLM_R_X15Y151_SLICE_X21Y151_CO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_C6 = CLBLM_R_X15Y153_SLICE_X21Y153_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_CIN = CLBLM_L_X16Y152_SLICE_X22Y152_COUT;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D6 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_CX = CLBLM_L_X16Y152_SLICE_X23Y152_CO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D1 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D2 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D3 = CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D4 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D5 = 1'b1;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_D6 = CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A1 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A2 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_DX = CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A4 = CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B2 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B3 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B4 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B5 = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B6 = CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C1 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C2 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C4 = CLBLM_R_X13Y131_SLICE_X18Y131_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C5 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C6 = CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D2 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A1 = CLBLM_R_X13Y138_SLICE_X19Y138_CQ;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A3 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B2 = CLBLM_R_X13Y137_SLICE_X19Y137_BQ;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B3 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B4 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B5 = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B6 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C1 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C2 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C3 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C4 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D1 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D2 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D3 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D4 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A1 = CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A3 = CLBLM_R_X13Y137_SLICE_X19Y137_AO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A4 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A6 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_AX = CLBLM_R_X13Y131_SLICE_X19Y131_CQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B1 = CLBLL_L_X26Y136_SLICE_X38Y136_BO5;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B3 = CLBLL_L_X26Y136_SLICE_X38Y136_BO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B4 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B6 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C1 = CLBLL_L_X26Y136_SLICE_X38Y136_BO5;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C2 = CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C3 = CLBLM_L_X12Y137_SLICE_X17Y137_BQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C6 = CLBLM_R_X13Y137_SLICE_X19Y137_BQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_CE = CLBLM_R_X13Y129_SLICE_X19Y129_AQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D2 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D3 = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D4 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D5 = CLBLM_R_X15Y137_SLICE_X21Y137_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D6 = CLBLM_R_X13Y134_SLICE_X19Y134_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A3 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_A6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_B6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C3 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_C6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B4 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B5 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D3 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X23Y154_D6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A1 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A3 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A4 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_A6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D5 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D6 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_AX = 1'b0;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B1 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B3 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B5 = CLBLL_L_X26Y133_SLICE_X38Y133_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B6 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C6 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_B5 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_BX = 1'b0;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A1 = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D4 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A2 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A3 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A4 = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A5 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_CX = 1'b0;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B1 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B2 = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A2 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A3 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A5 = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A6 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D1 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D2 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D3 = 1'b1;
  assign CLBLM_L_X16Y154_SLICE_X22Y154_D4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B1 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B3 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B4 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B6 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C1 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C2 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C3 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C1 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D1 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D2 = CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C2 = CLBLL_L_X26Y133_SLICE_X38Y133_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C4 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C5 = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C6 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D5 = CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D4 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A1 = CLBLM_R_X13Y138_SLICE_X19Y138_AQ;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A2 = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A4 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A5 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLL_L_X2Y144_SLICE_X0Y144_BQ;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B1 = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B2 = CLBLM_R_X13Y138_SLICE_X19Y138_BQ;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B4 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B5 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C2 = CLBLM_R_X13Y138_SLICE_X19Y138_CQ;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C3 = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C5 = CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C6 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X2Y144_SLICE_X0Y144_AQ;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D2 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A1 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A2 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A3 = CLBLM_R_X15Y137_SLICE_X21Y137_AQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A4 = CLBLM_R_X15Y138_SLICE_X21Y138_BQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A5 = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A6 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B1 = CLBLL_L_X26Y138_SLICE_X38Y138_AO5;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B2 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B3 = CLBLL_L_X26Y138_SLICE_X38Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B4 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B6 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C1 = CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C2 = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C3 = CLBLM_R_X13Y136_SLICE_X19Y136_BQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C4 = CLBLL_L_X26Y136_SLICE_X38Y136_BO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C6 = CLBLM_R_X13Y131_SLICE_X18Y131_BQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_CE = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D1 = CLBLM_L_X12Y136_SLICE_X17Y136_BQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D2 = CLBLM_R_X13Y131_SLICE_X18Y131_CQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D3 = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D4 = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D5 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D6 = CLBLL_L_X26Y138_SLICE_X38Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_D = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_D = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A2 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A3 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A4 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A5 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B2 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B3 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B4 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B5 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C1 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C4 = CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C5 = CLBLL_L_X26Y133_SLICE_X38Y133_DO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C6 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A1 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A3 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A4 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A6 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D4 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D6 = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D2 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A3 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A4 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B4 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B6 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C1 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C2 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C4 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C5 = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C6 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D1 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D2 = CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D4 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D6 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A1 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A2 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A3 = CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A4 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C4 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A5 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C5 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B1 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B2 = CLBLM_R_X13Y140_SLICE_X19Y140_BO5;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B3 = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B4 = CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C6 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B5 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B6 = CLBLM_R_X13Y139_SLICE_X19Y139_CO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C1 = CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B3 = CLBLL_L_X26Y133_SLICE_X38Y133_BO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C2 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C3 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C4 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C5 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B4 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C6 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D1 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D2 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D3 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D4 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D5 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D6 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_BI = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C1 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_CE = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C4 = CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D5 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D6 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C6 = CLBLL_L_X26Y133_SLICE_X38Y133_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_DI = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A5 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A1 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A2 = CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_AX = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D5 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D6 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C4 = CLBLM_R_X7Y138_SLICE_X8Y138_C_XOR;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C5 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A1 = CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A2 = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A3 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A5 = CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B1 = CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B3 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B4 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B5 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C1 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C2 = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C3 = CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C4 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C5 = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C6 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A1 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A3 = CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A4 = CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A5 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A6 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B1 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B2 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D5 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B3 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B4 = CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B5 = CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B6 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D3 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C1 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C2 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C3 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C4 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C5 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C6 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CE = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A1 = CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A3 = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A4 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D2 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D4 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D5 = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D6 = CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B2 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B5 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C1 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C3 = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C4 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C5 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CE = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D6 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D2 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D3 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A1 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A2 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A4 = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D3 = CLBLM_R_X15Y151_SLICE_X21Y151_AQ;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B1 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B5 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D4 = CLBLM_R_X15Y151_SLICE_X20Y151_AO5;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D5 = CLBLM_R_X15Y151_SLICE_X20Y151_BO5;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D6 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_AI = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_BI = CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_CE = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_CI = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D1 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D3 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_DI = 1'b0;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A3 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A4 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A5 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A6 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B1 = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B2 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B3 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B4 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B5 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B6 = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C1 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C3 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C5 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C6 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D1 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D2 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D3 = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D4 = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D5 = CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A1 = CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A3 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A4 = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A5 = CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A6 = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B1 = CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B2 = CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B3 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B4 = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B6 = CLBLM_R_X13Y137_SLICE_X18Y137_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D6 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C1 = CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C2 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A1 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C6 = CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_CE = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A3 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A4 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A5 = CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A6 = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C3 = CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_AX = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B1 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B2 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D2 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D3 = CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D4 = CLBLM_R_X13Y135_SLICE_X18Y135_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B3 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B4 = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B5 = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B6 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D5 = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C1 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C2 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C3 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C4 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C5 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C6 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A1 = CLBLM_R_X13Y138_SLICE_X19Y138_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A2 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A3 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A5 = LIOB33_X0Y187_IOB_X0Y188_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D1 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D2 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D3 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D4 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D5 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D6 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B2 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B3 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B4 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B5 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B6 = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C1 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C2 = CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C4 = CLBLM_L_X12Y137_SLICE_X16Y137_CO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C5 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C6 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D2 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D3 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D4 = CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A1 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_AX = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B1 = CLBLM_R_X15Y142_SLICE_X21Y142_DQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B2 = CLBLM_R_X15Y141_SLICE_X21Y141_BQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B3 = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B5 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B6 = CLBLM_L_X16Y142_SLICE_X22Y142_CQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_BX = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C1 = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C2 = CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C3 = CLBLM_R_X15Y143_SLICE_X20Y143_DO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C5 = CLBLM_R_X15Y139_SLICE_X20Y139_AO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C6 = CLBLM_R_X13Y141_SLICE_X19Y141_BO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_CE = CLBLM_L_X16Y141_SLICE_X22Y141_AO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_CX = CLBLM_R_X15Y139_SLICE_X21Y139_AO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D1 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D2 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D3 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D5 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D6 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A1 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A2 = CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A4 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A5 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A6 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B1 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B4 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B5 = CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B6 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C2 = CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C3 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C5 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C6 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D1 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D2 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D3 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D5 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A3 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B1 = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B3 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B4 = CLBLM_R_X7Y135_SLICE_X8Y135_AO5;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B5 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B6 = CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C1 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C2 = CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C3 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C4 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C5 = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C6 = CLBLM_R_X7Y134_SLICE_X9Y134_AO5;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D1 = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D3 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D4 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D5 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D6 = CLBLM_R_X7Y135_SLICE_X8Y135_AO5;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A1 = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A2 = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A3 = CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A4 = CLBLM_L_X8Y137_SLICE_X10Y137_AO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A6 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B1 = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B2 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B3 = CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B4 = CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B5 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B6 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A2 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A3 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_CE = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B1 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B2 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B3 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B4 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B5 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B6 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C1 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C2 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C3 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C5 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C6 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A2 = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D1 = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D2 = CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D3 = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D4 = CLBLM_R_X7Y134_SLICE_X8Y134_AO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D5 = CLBLL_L_X4Y135_SLICE_X5Y135_DO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D6 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B1 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B2 = CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B4 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B5 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C1 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C2 = CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C3 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C4 = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C5 = CLBLM_R_X15Y137_SLICE_X21Y137_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D1 = CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D2 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D3 = CLBLM_R_X15Y138_SLICE_X21Y138_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D4 = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D5 = CLBLM_R_X15Y144_SLICE_X20Y144_F7AMUX_O;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A2 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A3 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A4 = CLBLM_R_X13Y142_SLICE_X18Y142_BO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A5 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B1 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B2 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B3 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B5 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B6 = CLBLM_R_X11Y141_SLICE_X15Y141_AO5;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D1 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D2 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A1 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A2 = CLBLM_R_X15Y140_SLICE_X21Y140_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A3 = CLBLM_R_X15Y142_SLICE_X20Y142_BO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A4 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A5 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B1 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B2 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B3 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B4 = CLBLM_R_X15Y142_SLICE_X20Y142_AO5;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B5 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C1 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C3 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C4 = CLBLM_R_X15Y139_SLICE_X21Y139_AO5;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C5 = CLBLM_R_X15Y141_SLICE_X20Y141_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_CE = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D1 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D2 = CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D3 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D4 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D5 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A1 = CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A2 = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A4 = CLBLM_R_X11Y135_SLICE_X15Y135_AO5;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A5 = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A6 = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B1 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B4 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A3 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B5 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B6 = CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A4 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C2 = CLBLM_L_X10Y139_SLICE_X12Y139_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C1 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C3 = CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C5 = CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C6 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B1 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B3 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B4 = CLBLL_L_X4Y136_SLICE_X5Y136_DQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B5 = CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C1 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C2 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C3 = CLBLM_R_X15Y140_SLICE_X21Y140_AO5;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C4 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C5 = CLBLM_R_X15Y143_SLICE_X21Y143_AO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_CE = CLBLL_L_X2Y137_SLICE_X0Y137_BO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D2 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D3 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D4 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D2 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D3 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D4 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D5 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A1 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A2 = CLBLM_R_X15Y144_SLICE_X21Y144_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A4 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A5 = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_AX = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B1 = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B2 = CLBLM_R_X13Y131_SLICE_X18Y131_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B3 = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B4 = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B5 = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B6 = CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_BX = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C2 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C3 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C4 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D2 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D3 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D4 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D = LIOB33_X0Y181_IOB_X0Y181_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_D = LIOB33_X0Y197_IOB_X0Y197_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D = LIOB33_X0Y169_IOB_X0Y170_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A2 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A4 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A5 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_AX = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B2 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B4 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B5 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_BX = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C2 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C4 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C5 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_CE = CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_CX = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D2 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D4 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D5 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_DX = CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLL_L_X4Y135_SLICE_X4Y135_C5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A1 = CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A2 = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A3 = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A4 = CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A5 = CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A1 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A2 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A3 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A4 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A5 = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B4 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_AX = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B5 = CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B1 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_BX = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C5 = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C3 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C6 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_CE = CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CE = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D1 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_CX = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D2 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D4 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D5 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D4 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A1 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_DX = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A3 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A5 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B1 = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B2 = CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B3 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B4 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B5 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B6 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C1 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C2 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C3 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C5 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D2 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D3 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D4 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D5 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D6 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A1 = CLBLM_R_X13Y145_SLICE_X19Y145_BO5;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A2 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C2 = CLBLM_R_X13Y137_SLICE_X19Y137_AO5;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A6 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_AX = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B2 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B3 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B4 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B6 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C5 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C1 = CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C2 = CLBLM_R_X13Y144_SLICE_X18Y144_A_XOR;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C3 = CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C4 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C6 = CLBLL_L_X4Y137_SLICE_X5Y137_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C5 = CLBLM_R_X13Y145_SLICE_X18Y145_B_XOR;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B3 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D1 = CLBLM_R_X13Y144_SLICE_X18Y144_D_XOR;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B4 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D2 = CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D4 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D5 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D6 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A1 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A6 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_AX = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B1 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B2 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B4 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B6 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_BX = 1'b0;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C1 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C4 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C2 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_CX = 1'b0;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C3 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D1 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C4 = CLBLM_R_X13Y132_SLICE_X18Y132_BO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D6 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_DX = 1'b0;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D6 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C6 = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X15Y152_SLICE_X21Y152_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A1 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A2 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A4 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A5 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B1 = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B2 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B5 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B6 = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C1 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C2 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C3 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C4 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C5 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C6 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLL_L_X2Y135_SLICE_X1Y135_AQ;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_A5 = CLBLM_R_X15Y150_SLICE_X20Y150_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_AX = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D1 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D2 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D3 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D4 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D5 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D6 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_A6 = CLBLM_L_X16Y151_SLICE_X22Y151_A_XOR;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C2 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A1 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A1 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A2 = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A3 = CLBLL_L_X4Y137_SLICE_X5Y137_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A4 = CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A6 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A2 = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A3 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_BO5;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B1 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B2 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B3 = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B4 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B5 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B2 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B3 = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B4 = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C5 = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C6 = CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C2 = CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C3 = CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C5 = CLBLL_L_X4Y137_SLICE_X5Y137_BO5;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C6 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D2 = CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D6 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D1 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D3 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D4 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D5 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D6 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CE = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_C5 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_C6 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A1 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A2 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A4 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A5 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A6 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B1 = CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B2 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B3 = CLBLM_R_X13Y145_SLICE_X18Y145_C_XOR;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B4 = CLBLM_R_X13Y145_SLICE_X18Y145_A_XOR;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B5 = CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B6 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_D1 = CLBLM_L_X16Y133_SLICE_X23Y133_AQ;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C2 = CLBLM_R_X15Y146_SLICE_X20Y146_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C3 = CLBLM_R_X13Y144_SLICE_X19Y144_DO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C4 = CLBLM_R_X13Y145_SLICE_X19Y145_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C5 = CLBLM_R_X13Y148_SLICE_X18Y148_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C6 = CLBLM_R_X13Y146_SLICE_X19Y146_AO6;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_D5 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D4 = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_D6 = CLBLM_L_X16Y154_SLICE_X22Y154_A_CY;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D5 = CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D6 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A6 = 1'b1;
  assign CLBLM_R_X15Y152_SLICE_X20Y152_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_AX = 1'b0;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B6 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_BX = 1'b0;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C1 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C6 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_CIN = CLBLM_R_X13Y144_SLICE_X18Y144_COUT;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_CX = 1'b0;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D6 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_DX = 1'b0;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLL_L_X2Y135_SLICE_X1Y135_A5Q;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A1 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A2 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A3 = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A4 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A5 = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A1 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A2 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A3 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B1 = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B2 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B3 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B5 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A4 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_AX = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B4 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_BX = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C1 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C3 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C4 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D1 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D3 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D4 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D5 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D6 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A2 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A5 = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A4 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_AX = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B1 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B2 = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B3 = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B4 = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B5 = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B6 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_BX = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C1 = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C2 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C4 = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C5 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C6 = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D1 = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D2 = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D3 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D4 = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D6 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A3 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A5 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_A6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B1 = CLBLM_R_X13Y146_SLICE_X19Y146_DO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B2 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B3 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B4 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_B6 = CLBLM_R_X13Y146_SLICE_X19Y146_CO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C1 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C2 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C3 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C4 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_C6 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D2 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D4 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y146_SLICE_X19Y146_D6 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_AX = 1'b0;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_B6 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_BX = 1'b0;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C3 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_C6 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_CIN = CLBLM_R_X13Y145_SLICE_X18Y145_COUT;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_CX = 1'b0;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X4Y135_SLICE_X5Y135_A5Q;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D1 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D2 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D3 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D4 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D5 = 1'b1;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_D6 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_DX = 1'b0;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B3 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B4 = 1'b1;
  assign CLBLL_L_X2Y135_SLICE_X1Y135_B5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A1 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A2 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A3 = CLBLM_R_X11Y142_SLICE_X15Y142_F8MUX_O;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A4 = CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A5 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A6 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B1 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B2 = CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B3 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B4 = CLBLM_R_X11Y141_SLICE_X15Y141_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B5 = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B6 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C2 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C3 = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C4 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D1 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D3 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D4 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D5 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A1 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A3 = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A4 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A5 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A6 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B1 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B2 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B3 = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B4 = CLBLL_L_X4Y141_SLICE_X5Y141_CQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B5 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B6 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C1 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C2 = CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C3 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C4 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C5 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C6 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D1 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D2 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D3 = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D4 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D6 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A1 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A4 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A6 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B1 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B2 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B3 = CLBLM_R_X13Y148_SLICE_X19Y148_DO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B4 = CLBLM_R_X13Y147_SLICE_X19Y147_DO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B5 = CLBLM_R_X13Y147_SLICE_X19Y147_CO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B6 = CLBLM_R_X13Y148_SLICE_X19Y148_CO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C1 = CLBLM_R_X13Y147_SLICE_X19Y147_AO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C2 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C3 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C4 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C5 = CLBLM_L_X16Y152_SLICE_X23Y152_AO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C6 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D2 = CLBLM_R_X13Y146_SLICE_X19Y146_DO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D3 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D6 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_AX = 1'b0;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B6 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_BX = 1'b0;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C1 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C6 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_CIN = CLBLM_R_X13Y146_SLICE_X18Y146_COUT;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_CX = 1'b0;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D6 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_DX = 1'b0;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A2 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A3 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A4 = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C6 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_D1 = CLBLM_L_X16Y133_SLICE_X23Y133_BQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D6 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_D1 = CLBLM_L_X16Y133_SLICE_X22Y133_AQ;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A1 = CLBLL_L_X4Y141_SLICE_X5Y141_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A4 = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A5 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A6 = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_AX = CLBLM_R_X15Y142_SLICE_X20Y142_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B1 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B2 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B3 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A1 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A2 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_BX = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A6 = CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A3 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C3 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C6 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B4 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B5 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B6 = CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B1 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C2 = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C4 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C6 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D2 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_AX = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B1 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B2 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B3 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B4 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B5 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B6 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_BX = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C1 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C2 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C3 = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C4 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C6 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_CX = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D1 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D2 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D3 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D4 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D5 = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D6 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_DX = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A2 = CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A4 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A6 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B2 = CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B3 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B4 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B5 = CLBLM_R_X13Y148_SLICE_X19Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B6 = CLBLM_R_X13Y149_SLICE_X19Y149_AO5;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C2 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C3 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C4 = CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C5 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C6 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X2Y137_SLICE_X0Y137_AO6;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D = LIOB33_X0Y193_IOB_X0Y194_I;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D4 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D5 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D6 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D = LIOB33_X0Y193_IOB_X0Y193_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A1 = CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A2 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A3 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A5 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B1 = CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B2 = CLBLM_R_X15Y148_SLICE_X21Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B3 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B4 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B5 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B6 = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C1 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C2 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C3 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C4 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C5 = CLBLM_R_X13Y148_SLICE_X18Y148_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C6 = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D1 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D2 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D4 = CLBLM_L_X12Y144_SLICE_X16Y144_BO5;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D5 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D6 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A1 = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A2 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A4 = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A5 = CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A6 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_AX = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B1 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B3 = CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B5 = CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B6 = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C1 = CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C2 = CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C3 = CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C4 = CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C5 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D2 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D3 = CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D4 = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D5 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D6 = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A1 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A2 = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A4 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A5 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_AX = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B1 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B2 = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B4 = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B5 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_BX = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C1 = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C2 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C3 = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C4 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C5 = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A2 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A4 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B4 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B5 = CLBLM_R_X3Y141_SLICE_X3Y141_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B6 = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_AX = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_CX = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B1 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C2 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C3 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C4 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C5 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D2 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D3 = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D5 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_DX = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D1 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D3 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A2 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A3 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A4 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A6 = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_AX = CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B1 = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B3 = CLBLM_R_X3Y141_SLICE_X3Y141_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B4 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B6 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_BX = CLBLM_L_X10Y144_SLICE_X13Y144_DO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C1 = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C2 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C3 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C4 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C5 = CLBLM_R_X3Y141_SLICE_X3Y141_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C6 = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CIN = CLBLM_L_X10Y144_SLICE_X12Y144_COUT;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CX = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D4 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D5 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D6 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_DX = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B4 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B5 = CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B6 = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X2Y137_SLICE_X1Y137_AO6;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLL_L_X2Y137_SLICE_X0Y137_AO5;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A1 = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A2 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A3 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B4 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B5 = CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B6 = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C5 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B1 = CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C6 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A1 = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A2 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A3 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A4 = CLBLM_R_X15Y153_SLICE_X21Y153_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C4 = CLBLM_L_X12Y131_SLICE_X16Y131_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B1 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B2 = CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B3 = CLBLM_R_X13Y148_SLICE_X18Y148_AO5;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C6 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C1 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A3 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A4 = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A6 = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C2 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A1 = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A2 = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A3 = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A4 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A6 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B1 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AX = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B2 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B1 = CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B3 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B4 = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B6 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B5 = CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C1 = CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C2 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C4 = CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C5 = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C6 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CE = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D3 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D4 = CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D5 = CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D6 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B1 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B2 = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B6 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A1 = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A2 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A3 = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A4 = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A5 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_AX = CLBLM_R_X3Y141_SLICE_X3Y141_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B1 = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B2 = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B3 = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B4 = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B5 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_BX = CLBLM_R_X3Y141_SLICE_X3Y141_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C1 = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C2 = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C3 = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C4 = CLBLM_R_X3Y141_SLICE_X3Y141_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C5 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CIN = CLBLL_L_X4Y141_SLICE_X5Y141_COUT;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A2 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A3 = CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A4 = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A5 = CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CX = CLBLM_R_X3Y141_SLICE_X3Y141_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A6 = CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B2 = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B3 = CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B4 = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B6 = CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D3 = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D4 = CLBLM_R_X3Y141_SLICE_X3Y141_DQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C2 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C3 = CLBLM_L_X12Y143_SLICE_X16Y143_BO5;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C4 = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C5 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C6 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_DX = CLBLM_R_X3Y141_SLICE_X3Y141_DQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C1 = CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_CE = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D2 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D4 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D6 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A1 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A3 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A4 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A5 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A6 = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_AX = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B1 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B3 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B4 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B6 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_BX = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C2 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C4 = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C6 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = CLBLM_L_X16Y133_SLICE_X22Y133_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CIN = CLBLM_L_X10Y145_SLICE_X12Y145_COUT;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CX = CLBLM_L_X10Y147_SLICE_X13Y147_DO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D2 = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D3 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D4 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D6 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X2Y137_SLICE_X1Y137_AO5;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X2Y137_SLICE_X1Y137_BO6;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_DX = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A1 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A2 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A3 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A4 = CLBLM_R_X15Y151_SLICE_X20Y151_CO5;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A6 = CLBLM_R_X13Y150_SLICE_X19Y150_CO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_AX = CLBLM_R_X15Y150_SLICE_X20Y150_DO5;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B1 = CLBLM_R_X13Y150_SLICE_X19Y150_DO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B5 = CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B6 = CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C2 = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C4 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C5 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C6 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D1 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D2 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D5 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D6 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A1 = CLBLM_R_X15Y150_SLICE_X20Y150_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D6 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A2 = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A3 = CLBLM_R_X15Y150_SLICE_X21Y150_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C5 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B6 = CLBLM_R_X5Y149_SLICE_X6Y149_AO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B1 = CLBLM_R_X13Y150_SLICE_X18Y150_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B3 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_DX = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C3 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C4 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C6 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D2 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A2 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A1 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A2 = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A3 = CLBLM_R_X15Y148_SLICE_X21Y148_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A4 = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A5 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A6 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A3 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A4 = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A5 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B1 = CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B2 = CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B4 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B5 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B6 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B2 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B4 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C1 = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C2 = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C4 = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C5 = CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C6 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C1 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C2 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C3 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C4 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C5 = CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C6 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CE = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D1 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D2 = CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D3 = CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D4 = CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D6 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D1 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D2 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D3 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D4 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D6 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A2 = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A3 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A6 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_AX = 1'b0;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B6 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_BX = 1'b0;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C6 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CIN = CLBLL_L_X4Y142_SLICE_X5Y142_COUT;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A1 = CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A2 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A3 = CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A4 = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CX = 1'b0;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D6 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B5 = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B6 = CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_DX = 1'b0;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B2 = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B3 = CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B4 = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C3 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C4 = CLBLM_L_X10Y147_SLICE_X13Y147_AO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C5 = CLBLM_L_X12Y146_SLICE_X17Y146_F7AMUX_O;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C6 = CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C1 = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C2 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D5 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D2 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D3 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D4 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D5 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A2 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A4 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A5 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A6 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y139_SLICE_X1Y139_DO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X2Y137_SLICE_X1Y137_BO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_AX = CLBLM_R_X11Y147_SLICE_X14Y147_DO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B1 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B2 = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B3 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B4 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B6 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_BX = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C2 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C4 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C5 = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C6 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CIN = CLBLM_L_X10Y146_SLICE_X12Y146_COUT;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CX = 1'b0;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D2 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D3 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D4 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D5 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_DX = 1'b0;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A1 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A4 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A5 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A6 = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B1 = CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B2 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B3 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B4 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B5 = CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B6 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A1 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A2 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A4 = CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A5 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A6 = CLBLM_R_X3Y142_SLICE_X3Y142_DQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A1 = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A2 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A3 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B3 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B4 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B5 = CLBLL_L_X2Y157_SLICE_X0Y157_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A5 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A6 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C1 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C2 = CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C3 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C4 = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C6 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B4 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B5 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B6 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C1 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C4 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D2 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D3 = CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D4 = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D6 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D1 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D4 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D6 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A4 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_AX = 1'b0;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B2 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B5 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_BX = 1'b0;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C6 = CLBLM_R_X3Y143_SLICE_X3Y143_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CIN = CLBLL_L_X4Y143_SLICE_X5Y143_COUT;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CX = 1'b0;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A1 = CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D6 = CLBLM_R_X3Y143_SLICE_X3Y143_DQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A2 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A3 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_DX = 1'b0;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A4 = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B6 = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B5 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C4 = CLBLM_R_X13Y147_SLICE_X18Y147_B_XOR;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C5 = CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C6 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C2 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X2Y139_SLICE_X1Y139_DO5;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLL_L_X2Y139_SLICE_X1Y139_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D4 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A1 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A2 = CLBLM_R_X13Y147_SLICE_X18Y147_C_XOR;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A3 = CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A4 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B2 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B5 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B6 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C1 = CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C2 = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C3 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C4 = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C6 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D4 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D6 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = CLBLM_L_X16Y134_SLICE_X23Y134_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A1 = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A6 = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B6 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C6 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = CLBLM_L_X16Y133_SLICE_X23Y133_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A3 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A4 = CLBLL_L_X2Y156_SLICE_X0Y156_BO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A5 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A1 = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B1 = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B2 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B4 = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B5 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B6 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A2 = CLBLM_R_X13Y144_SLICE_X19Y144_F7AMUX_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A3 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A4 = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C1 = CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C2 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C3 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B1 = CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B2 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C1 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C2 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C4 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D1 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D2 = CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D3 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D6 = CLBLL_L_X4Y142_SLICE_X5Y142_DQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C6 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D1 = CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D2 = CLBLM_R_X5Y129_SLICE_X6Y129_DQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D4 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D5 = CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D6 = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C1 = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A1 = CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A2 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A3 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A4 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A5 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C2 = CLBLM_L_X16Y137_SLICE_X22Y137_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B1 = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B3 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B4 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B5 = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B6 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C1 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C2 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C3 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C4 = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C5 = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C6 = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C3 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLL_L_X2Y139_SLICE_X1Y139_BO6;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X2Y139_SLICE_X1Y139_AO5;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D2 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D4 = CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A1 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A2 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A4 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A5 = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A6 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_BO5;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D6 = CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B1 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B2 = CLBLM_L_X10Y150_SLICE_X13Y150_AO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B3 = CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B4 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B5 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B6 = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C4 = CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C1 = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C4 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C5 = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C6 = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D2 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D3 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D4 = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D5 = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D6 = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A2 = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A4 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A6 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B2 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B3 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B4 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C6 = CLBLM_L_X16Y137_SLICE_X22Y137_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C2 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C3 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C4 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D2 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D3 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D4 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A2 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A3 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A4 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A5 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A6 = CLBLM_L_X10Y135_SLICE_X12Y135_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B1 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B2 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B3 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B5 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B6 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C2 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A1 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A5 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D2 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B3 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B5 = CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B6 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A2 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A3 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C2 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C3 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C4 = CLBLL_L_X2Y155_SLICE_X0Y155_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A6 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B1 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B2 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B3 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B4 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C1 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C4 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C6 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D2 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A1 = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A2 = CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A3 = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A6 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X2Y139_SLICE_X1Y139_CO6;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X2Y139_SLICE_X1Y139_BO5;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B3 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C3 = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A1 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A2 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A5 = CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B2 = CLBLM_R_X15Y150_SLICE_X21Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B4 = CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B5 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B6 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C3 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D3 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A3 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B3 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C3 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D3 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B1 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B2 = CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B5 = CLBLM_R_X15Y145_SLICE_X20Y145_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_BX = CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B3 = CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C1 = CLBLM_R_X15Y142_SLICE_X20Y142_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B4 = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C2 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C3 = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B6 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A2 = CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A3 = CLBLM_L_X16Y136_SLICE_X22Y136_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A4 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A5 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B1 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B2 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B3 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B4 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B5 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B6 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B3 = CLBLM_R_X15Y137_SLICE_X21Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B4 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C1 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C3 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C4 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C6 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B5 = CLBLM_R_X13Y137_SLICE_X18Y137_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A2 = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A3 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A4 = CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C4 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A6 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C5 = CLBLM_L_X12Y130_SLICE_X16Y130_CQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B1 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B2 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B3 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B4 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C6 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B6 = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A1 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_CE = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C2 = CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C3 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C5 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C6 = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A3 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A4 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A5 = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A6 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D5 = CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D6 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B4 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C1 = CLBLL_L_X4Y136_SLICE_X5Y136_DQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C2 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C4 = CLBLM_R_X5Y141_SLICE_X7Y141_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C5 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C6 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D5 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D6 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C5 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D2 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D4 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D5 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D6 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A1 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A4 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A6 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B1 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B3 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B4 = CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B6 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = CLBLM_L_X16Y134_SLICE_X22Y134_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C1 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C2 = CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C3 = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C4 = CLBLL_L_X4Y147_SLICE_X5Y147_AO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C6 = CLBLL_L_X4Y149_SLICE_X5Y149_AO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D3 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D5 = CLBLM_R_X5Y148_SLICE_X7Y148_BO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = CLBLM_L_X16Y135_SLICE_X22Y135_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A2 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A4 = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A6 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B3 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B4 = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B6 = CLBLM_R_X15Y151_SLICE_X20Y151_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D6 = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D6 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_A1 = CLBLL_L_X2Y138_SLICE_X0Y138_B_XOR;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A1 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A2 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A3 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A4 = CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A5 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A6 = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_AX = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B1 = CLBLM_R_X15Y145_SLICE_X20Y145_F7AMUX_O;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B2 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B3 = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B5 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B6 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D4 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C1 = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C2 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C3 = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B2 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C4 = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A6 = 1'b1;
  assign CLBLL_L_X2Y137_SLICE_X0Y137_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y116_SLICE_X0Y116_B1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B3 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B5 = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D1 = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C4 = CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C5 = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D4 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A1 = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A2 = CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A4 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A5 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D4 = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B2 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B3 = CLBLM_L_X12Y130_SLICE_X16Y130_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B4 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B5 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B6 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C2 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C3 = CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C4 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C5 = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C6 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D1 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D3 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D4 = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D5 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D6 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A1 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A3 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A4 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B1 = CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B2 = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B3 = CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B4 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B5 = CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B6 = CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C1 = CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C2 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C4 = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C5 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_CE = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D1 = CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D2 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D5 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A1 = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A2 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A3 = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A4 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A5 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B2 = CLBLM_L_X8Y134_SLICE_X10Y134_F8MUX_O;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B3 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B4 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B5 = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B6 = CLBLM_R_X11Y137_SLICE_X14Y137_F8MUX_O;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A2 = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A3 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A5 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C1 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C2 = CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C3 = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B3 = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B4 = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B5 = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B6 = CLBLL_L_X4Y149_SLICE_X4Y149_AO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D2 = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C6 = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D3 = CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A1 = CLBLM_L_X12Y151_SLICE_X17Y151_F8MUX_O;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A2 = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A3 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A4 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A5 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D3 = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D5 = CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B1 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B2 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B4 = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B5 = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B6 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C1 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C2 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C4 = CLBLM_R_X5Y137_SLICE_X7Y137_BO5;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C5 = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C6 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D1 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D2 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D3 = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A5 = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D6 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B1 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B3 = CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B4 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B5 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B6 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C2 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C4 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C5 = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C6 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D1 = CLBLM_R_X5Y151_SLICE_X6Y151_BO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D2 = CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D6 = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D6 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = CLBLM_L_X16Y135_SLICE_X22Y135_BQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = CLBLM_L_X16Y135_SLICE_X23Y135_AQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X2Y144_SLICE_X0Y144_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A1 = CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A2 = CLBLM_R_X15Y140_SLICE_X21Y140_AO5;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A4 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A5 = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B2 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B3 = CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B4 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B5 = CLBLL_L_X4Y138_SLICE_X5Y138_AO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A2 = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A3 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A4 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A5 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B6 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_AX = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B2 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B5 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B6 = CLBLM_R_X3Y140_SLICE_X2Y140_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C4 = CLBLL_L_X4Y138_SLICE_X5Y138_AO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_BX = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C2 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C3 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C4 = CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C5 = CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C6 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_CE = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D3 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D4 = CLBLM_L_X16Y137_SLICE_X22Y137_BO5;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D5 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_CX = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A1 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D1 = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D2 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D3 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D4 = CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D5 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D6 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A3 = CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A4 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A5 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A6 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_AX = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B1 = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B2 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B4 = CLBLL_L_X4Y137_SLICE_X5Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B5 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B6 = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C1 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C2 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C3 = CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C4 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C5 = CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C6 = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A1 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A4 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D2 = CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D3 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B1 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B2 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B3 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B6 = CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D1 = CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLL_L_X2Y145_SLICE_X0Y145_AQ;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X2Y144_SLICE_X0Y144_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A1 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A2 = CLBLM_R_X7Y138_SLICE_X8Y138_D_XOR;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A3 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A4 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A5 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A6 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A1 = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A2 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A3 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A4 = CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A5 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A6 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B1 = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B2 = CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_AX = CLBLL_L_X4Y151_SLICE_X4Y151_DO5;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B3 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B1 = CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B2 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B3 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B4 = CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B5 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B6 = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_BX = CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C1 = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C2 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C1 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C2 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C3 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C4 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C5 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C6 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D1 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D3 = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D4 = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D5 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D2 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D3 = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D4 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D5 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A1 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_SR = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A3 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A5 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_AX = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B2 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B3 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B4 = CLBLM_R_X15Y144_SLICE_X21Y144_AO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B5 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B6 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_BX = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C1 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C2 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C3 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C4 = CLBLM_R_X15Y144_SLICE_X20Y144_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C5 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C6 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_B5 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A1 = CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A2 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A3 = CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A4 = CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A5 = CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A6 = CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_CX = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D1 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D2 = CLBLM_R_X15Y144_SLICE_X21Y144_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B1 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B5 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D3 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D4 = CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D5 = CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C5 = CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X15Y150_SLICE_X20Y150_B6 = CLBLM_R_X15Y150_SLICE_X20Y150_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_COUT = CLBLL_L_X2Y138_SLICE_X0Y138_D_CY;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_COUT = CLBLL_L_X2Y139_SLICE_X0Y139_D_CY;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_COUT = CLBLL_L_X2Y140_SLICE_X0Y140_D_CY;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_COUT = CLBLL_L_X2Y140_SLICE_X1Y140_D_CY;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_COUT = CLBLL_L_X2Y141_SLICE_X1Y141_D_CY;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_COUT = CLBLL_L_X2Y142_SLICE_X1Y142_D_CY;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_COUT = CLBLL_L_X4Y141_SLICE_X5Y141_D_CY;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_COUT = CLBLL_L_X4Y142_SLICE_X5Y142_D_CY;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_COUT = CLBLL_L_X4Y143_SLICE_X5Y143_D_CY;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_COUT = CLBLM_L_X10Y144_SLICE_X12Y144_D_CY;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_COUT = CLBLM_L_X10Y145_SLICE_X12Y145_D_CY;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_COUT = CLBLM_L_X10Y146_SLICE_X12Y146_D_CY;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_COUT = CLBLM_L_X12Y147_SLICE_X16Y147_D_CY;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_COUT = CLBLM_L_X12Y147_SLICE_X17Y147_D_CY;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_COUT = CLBLM_L_X12Y148_SLICE_X16Y148_D_CY;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_COUT = CLBLM_L_X12Y148_SLICE_X17Y148_D_CY;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_COUT = CLBLM_L_X12Y149_SLICE_X17Y149_D_CY;
  assign CLBLM_L_X16Y150_SLICE_X22Y150_COUT = CLBLM_L_X16Y150_SLICE_X22Y150_D_CY;
  assign CLBLM_L_X16Y152_SLICE_X22Y152_COUT = CLBLM_L_X16Y152_SLICE_X22Y152_D_CY;
  assign CLBLM_L_X16Y153_SLICE_X22Y153_COUT = CLBLM_L_X16Y153_SLICE_X22Y153_D_CY;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_COUT = CLBLM_R_X3Y140_SLICE_X3Y140_D_CY;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_COUT = CLBLM_R_X3Y141_SLICE_X3Y141_D_CY;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_COUT = CLBLM_R_X3Y142_SLICE_X3Y142_D_CY;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_COUT = CLBLM_R_X5Y128_SLICE_X7Y128_D_CY;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_COUT = CLBLM_R_X5Y129_SLICE_X7Y129_D_CY;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_COUT = CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_COUT = CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_COUT = CLBLM_R_X5Y131_SLICE_X6Y131_D_CY;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_COUT = CLBLM_R_X5Y132_SLICE_X6Y132_D_CY;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_COUT = CLBLM_R_X5Y142_SLICE_X6Y142_D_CY;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_COUT = CLBLM_R_X5Y143_SLICE_X6Y143_D_CY;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_COUT = CLBLM_R_X7Y138_SLICE_X8Y138_D_CY;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_COUT = CLBLM_R_X11Y130_SLICE_X14Y130_D_CY;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_COUT = CLBLM_R_X11Y130_SLICE_X15Y130_D_CY;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_COUT = CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_COUT = CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_COUT = CLBLM_R_X11Y132_SLICE_X14Y132_D_CY;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_COUT = CLBLM_R_X11Y132_SLICE_X15Y132_D_CY;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_COUT = CLBLM_R_X13Y144_SLICE_X18Y144_D_CY;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_COUT = CLBLM_R_X13Y145_SLICE_X18Y145_D_CY;
  assign CLBLM_R_X13Y146_SLICE_X18Y146_COUT = CLBLM_R_X13Y146_SLICE_X18Y146_D_CY;
  assign CLBLM_R_X15Y134_SLICE_X20Y134_COUT = CLBLM_R_X15Y134_SLICE_X20Y134_D_CY;
  assign CLBLM_R_X15Y135_SLICE_X20Y135_COUT = CLBLM_R_X15Y135_SLICE_X20Y135_D_CY;
  assign CLBLM_R_X15Y136_SLICE_X20Y136_COUT = CLBLM_R_X15Y136_SLICE_X20Y136_D_CY;
endmodule
