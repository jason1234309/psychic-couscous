module top(
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output RIOB33_SING_X105Y149_IOB_X1Y149_OPAD,
  output RIOB33_X105Y115_IOB_X1Y115_OPAD,
  output RIOB33_X105Y115_IOB_X1Y116_OPAD,
  output RIOB33_X105Y117_IOB_X1Y117_OPAD,
  output RIOB33_X105Y117_IOB_X1Y118_OPAD,
  output RIOB33_X105Y119_IOB_X1Y119_OPAD,
  output RIOB33_X105Y119_IOB_X1Y120_OPAD,
  output RIOB33_X105Y121_IOB_X1Y121_OPAD,
  output RIOB33_X105Y121_IOB_X1Y122_OPAD,
  output RIOB33_X105Y123_IOB_X1Y123_OPAD,
  output RIOB33_X105Y123_IOB_X1Y124_OPAD,
  output RIOB33_X105Y125_IOB_X1Y125_OPAD,
  output RIOB33_X105Y125_IOB_X1Y126_OPAD,
  output RIOB33_X105Y127_IOB_X1Y127_OPAD,
  output RIOB33_X105Y129_IOB_X1Y129_OPAD,
  output RIOB33_X105Y129_IOB_X1Y130_OPAD,
  output RIOB33_X105Y131_IOB_X1Y131_OPAD,
  output RIOB33_X105Y131_IOB_X1Y132_OPAD,
  output RIOB33_X105Y133_IOB_X1Y133_OPAD,
  output RIOB33_X105Y133_IOB_X1Y134_OPAD,
  output RIOB33_X105Y135_IOB_X1Y135_OPAD,
  output RIOB33_X105Y135_IOB_X1Y136_OPAD,
  output RIOB33_X105Y137_IOB_X1Y137_OPAD,
  output RIOB33_X105Y137_IOB_X1Y138_OPAD,
  output RIOB33_X105Y139_IOB_X1Y139_OPAD,
  output RIOB33_X105Y139_IOB_X1Y140_OPAD,
  output RIOB33_X105Y141_IOB_X1Y141_OPAD,
  output RIOB33_X105Y141_IOB_X1Y142_OPAD,
  output RIOB33_X105Y143_IOB_X1Y143_OPAD,
  output RIOB33_X105Y143_IOB_X1Y144_OPAD,
  output RIOB33_X105Y145_IOB_X1Y145_OPAD,
  output RIOB33_X105Y145_IOB_X1Y146_OPAD,
  output RIOB33_X105Y147_IOB_X1Y147_OPAD,
  output RIOB33_X105Y147_IOB_X1Y148_OPAD
  );
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A1;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A2;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A3;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A4;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A5Q;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_AMUX;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_AO5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_AO6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_AQ;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A_CY;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_A_XOR;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_B;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_B1;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_B2;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_B3;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_B4;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_B5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_B6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_BO5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_BO6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_BQ;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_B_CY;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_B_XOR;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_C;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_C1;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_C2;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_C3;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_C4;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_C5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_C6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_CLK;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_CO5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_CO6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_CQ;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_C_CY;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_C_XOR;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_D;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_D1;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_D2;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_D3;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_D4;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_D5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_D6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_DO5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_DO6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_D_CY;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_D_XOR;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X160Y107_SR;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_A;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_A1;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_A2;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_A3;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_A4;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_A5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_A6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_AO5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_AO6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_A_CY;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_A_XOR;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_B;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_B1;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_B2;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_B3;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_B4;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_B5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_B6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_BO5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_BO6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_B_CY;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_B_XOR;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_C;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_C1;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_C2;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_C3;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_C4;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_C5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_C6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_CO5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_CO6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_C_CY;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_C_XOR;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_D;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_D1;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_D2;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_D3;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_D4;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_D5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_D6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_DO5;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_DO6;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_D_CY;
  wire [0:0] CLBLL_L_X102Y107_SLICE_X161Y107_D_XOR;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_A;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_A1;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_A2;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_A3;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_A4;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_A5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_A6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_AO5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_AO6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_A_CY;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_A_XOR;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_B;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_B1;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_B2;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_B3;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_B4;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_B5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_B6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_BO5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_BO6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_B_CY;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_B_XOR;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_C;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_C1;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_C2;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_C3;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_C4;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_C5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_C6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_CO5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_CO6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_C_CY;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_C_XOR;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_D;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_D1;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_D2;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_D3;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_D4;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_D5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_D6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_DO5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_DO6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_D_CY;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X160Y108_D_XOR;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_A;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_A1;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_A2;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_A3;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_A4;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_A5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_A6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_AO5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_AO6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_AQ;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_A_CY;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_A_XOR;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B1;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B2;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B3;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B4;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B5Q;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_BMUX;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_BO5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_BO6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_BQ;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B_CY;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_B_XOR;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_C;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_C1;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_C2;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_C3;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_C4;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_C5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_C6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_CLK;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_CO5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_CO6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_C_CY;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_C_XOR;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_D;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_D1;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_D2;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_D3;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_D4;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_D5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_D6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_DO5;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_DO6;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_D_CY;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_D_XOR;
  wire [0:0] CLBLL_L_X102Y108_SLICE_X161Y108_SR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A1;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A2;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A3;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A4;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A5Q;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_AMUX;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_AO5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_AO6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_AQ;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A_CY;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_A_XOR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B1;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B2;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B3;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B4;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B5Q;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_BMUX;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_BO5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_BO6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_BQ;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B_CY;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_B_XOR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C1;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C2;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C3;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C4;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C5Q;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_CLK;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_CMUX;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_CO5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_CO6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_CQ;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C_CY;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_C_XOR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_D;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_D1;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_D2;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_D3;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_D4;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_D5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_D6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_DO5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_DO6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_D_CY;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_D_XOR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X160Y109_SR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_A;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_A1;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_A2;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_A3;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_A4;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_A5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_A6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_AMUX;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_AO5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_AO6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_AQ;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_A_CY;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_A_XOR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B1;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B2;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B3;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B4;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B5Q;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_BMUX;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_BO5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_BO6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_BQ;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B_CY;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_B_XOR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_C;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_C1;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_C2;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_C3;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_C4;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_C5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_C6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_CLK;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_CMUX;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_CO5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_CO6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_CQ;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_C_CY;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_C_XOR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_D;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_D1;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_D2;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_D3;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_D4;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_D5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_D6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_DO5;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_DO6;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_DQ;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_DX;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_D_CY;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_D_XOR;
  wire [0:0] CLBLL_L_X102Y109_SLICE_X161Y109_SR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A1;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A2;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A3;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A4;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A5Q;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_AMUX;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_AO5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_AO6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_AQ;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A_CY;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_A_XOR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B1;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B2;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B3;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B4;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B5Q;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_BMUX;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_BO5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_BO6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_BQ;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B_CY;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_B_XOR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C1;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C2;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C3;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C4;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C5Q;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_CLK;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_CMUX;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_CO5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_CO6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_CQ;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C_CY;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_C_XOR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D1;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D2;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D3;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D4;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D5Q;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_DMUX;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_DO5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_DO6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_DQ;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D_CY;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_D_XOR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X160Y110_SR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A1;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A2;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A3;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A4;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A5Q;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_AMUX;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_AO5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_AO6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_AQ;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A_CY;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_A_XOR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B1;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B2;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B3;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B4;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B5Q;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_BMUX;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_BO5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_BO6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_BQ;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B_CY;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_B_XOR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_C;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_C1;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_C2;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_C3;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_C4;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_C5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_C6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_CLK;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_CO5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_CO6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_CQ;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_CX;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_C_CY;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_C_XOR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_D;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_D1;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_D2;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_D3;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_D4;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_D5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_D6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_DO5;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_DO6;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_D_CY;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_D_XOR;
  wire [0:0] CLBLL_L_X102Y110_SLICE_X161Y110_SR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A5Q;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_AMUX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_AO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_AO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_AQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_AX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_A_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B5Q;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_BMUX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_BO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_BO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_BQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_BX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_B_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C5Q;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CLK;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CMUX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_CX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_C_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_DO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_DO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_DQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_DX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_D_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X160Y111_SR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_AO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_AO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_AQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_AX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_A_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_BO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_BO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_BQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_BX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_B_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CLK;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_CX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_C_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D1;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D2;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D3;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D4;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_DO5;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_DO6;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_DQ;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_DX;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D_CY;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_D_XOR;
  wire [0:0] CLBLL_L_X102Y111_SLICE_X161Y111_SR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A5Q;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_AMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_AO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_AO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_AX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_A_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B5Q;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_BMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_BO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_BO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_BX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_B_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C5Q;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CLK;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_CX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_C_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_DO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_DO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_DQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_DX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_D_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X160Y112_SR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A5Q;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_AMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_AO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_AO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_AQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_AX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_A_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B5Q;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_BMUX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_BO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_BO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_BX;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_B_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_CLK;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_CO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_CO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_C_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D1;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D2;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D3;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D4;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_DO5;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_DO6;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D_CY;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_D_XOR;
  wire [0:0] CLBLL_L_X102Y112_SLICE_X161Y112_SR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_AO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_AO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_A_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_BO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_BO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_B_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_CO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_CO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_C_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_DO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_DO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X160Y113_D_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_AO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_AO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_A_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_BO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_BO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_B_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_CLK;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_CO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_CO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_C_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D1;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D2;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D3;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D4;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_DO5;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_DO6;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D_CY;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_D_XOR;
  wire [0:0] CLBLL_L_X102Y113_SLICE_X161Y113_SR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_AO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_AO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_A_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_BO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_BO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_B_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_CO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_CO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_C_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_DO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_DO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X160Y114_D_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_AO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_AO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_AQ;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_A_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_BO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_BO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_B_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_CLK;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_CO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_CO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_C_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D1;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D2;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D3;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D4;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_DO5;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_DO6;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D_CY;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_D_XOR;
  wire [0:0] CLBLL_L_X102Y114_SLICE_X161Y114_SR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_AO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_AO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_AQ;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_A_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_BO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_BO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_B_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_CLK;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_CO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_CO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_C_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_DO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_DO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_D_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X160Y115_SR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_AMUX;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_AO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_AO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_AQ;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_AX;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_A_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_BO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_BO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_BQ;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_B_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_CLK;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_CO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_CO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_CQ;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_C_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D1;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D2;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D3;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D4;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_DO5;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_DO6;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D_CY;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_D_XOR;
  wire [0:0] CLBLL_L_X102Y115_SLICE_X161Y115_SR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A5Q;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_AMUX;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_AO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_AO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_AQ;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_A_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B5Q;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_BMUX;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_BO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_BO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_BQ;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_B_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_CLK;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_CMUX;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_CO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_CO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_C_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_DO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_DO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_D_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X162Y108_SR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AQ;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_AX;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_A_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_BO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_BO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_B_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_CLK;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_CO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_CO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_C_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D1;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D2;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D3;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D4;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_DO5;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_DO6;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D_CY;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_D_XOR;
  wire [0:0] CLBLM_R_X103Y108_SLICE_X163Y108_SR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A1;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A2;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A3;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A4;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A5Q;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_AMUX;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_AO5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_AO6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_AQ;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A_CY;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_A_XOR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B1;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B2;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B3;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B4;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B5Q;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_BMUX;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_BO5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_BO6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_BQ;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B_CY;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_B_XOR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_C;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_C1;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_C2;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_C3;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_C4;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_C5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_C6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_CLK;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_CMUX;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_CO5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_CO6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_CQ;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_C_CY;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_C_XOR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_D;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_D1;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_D2;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_D3;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_D4;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_D5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_D6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_DO5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_DO6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_D_CY;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_D_XOR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X162Y109_SR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_A;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_A1;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_A2;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_A3;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_A4;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_A5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_A6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_AMUX;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_AO5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_AO6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_AQ;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_A_CY;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_A_XOR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B1;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B2;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B3;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B4;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B5Q;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_BMUX;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_BO5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_BO6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_BQ;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B_CY;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_B_XOR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_C;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_C1;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_C2;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_C3;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_C4;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_C5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_C6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_CLK;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_CO5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_CO6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_CQ;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_C_CY;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_C_XOR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_D;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_D1;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_D2;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_D3;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_D4;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_D5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_D6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_DO5;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_DO6;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_D_CY;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_D_XOR;
  wire [0:0] CLBLM_R_X103Y109_SLICE_X163Y109_SR;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A1;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A2;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A3;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A4;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A5Q;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_AMUX;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_AO5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_AO6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_AQ;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A_CY;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_A_XOR;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B1;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B2;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B3;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B4;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B5Q;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_BMUX;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_BO5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_BO6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_BQ;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B_CY;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_B_XOR;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C1;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C2;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C3;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C4;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C5Q;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_CLK;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_CMUX;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_CO5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_CO6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_CQ;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C_CY;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_C_XOR;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D1;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D2;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D3;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D4;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D5Q;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_DMUX;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_DO5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_DO6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_DQ;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D_CY;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_D_XOR;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X162Y110_SR;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_A;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_A1;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_A2;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_A3;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_A4;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_A5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_A6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_AO5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_AO6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_A_CY;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_A_XOR;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_B;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_B1;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_B2;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_B3;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_B4;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_B5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_B6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_BO5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_BO6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_B_CY;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_B_XOR;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_C;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_C1;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_C2;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_C3;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_C4;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_C5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_C6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_CO5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_CO6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_C_CY;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_C_XOR;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_D;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_D1;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_D2;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_D3;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_D4;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_D5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_D6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_DO5;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_DO6;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_D_CY;
  wire [0:0] CLBLM_R_X103Y110_SLICE_X163Y110_D_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A5Q;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_AMUX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_AO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_AO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_AQ;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_A_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B5Q;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_BMUX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_BO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_BO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_BQ;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_B_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_CLK;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_CO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_CO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_C_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_DO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_DO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_D_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X162Y111_SR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_AO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_AO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_AQ;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_AX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_A_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_BO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_BO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_BQ;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_BX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_B_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_CLK;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_CO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_CO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_CQ;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_CX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_C_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D1;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D2;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D3;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D4;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_DO5;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_DO6;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_DQ;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_DX;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D_CY;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_D_XOR;
  wire [0:0] CLBLM_R_X103Y111_SLICE_X163Y111_SR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_AMUX;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_AO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_AO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_AQ;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_A_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_BO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_BO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_B_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_CLK;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_CO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_CO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_C_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_DO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_DO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_D_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X162Y112_SR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_AO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_AO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_A_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_BO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_BO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_B_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_CO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_CO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_C_XOR;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D1;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D2;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D3;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D4;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_DO5;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_DO6;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D_CY;
  wire [0:0] CLBLM_R_X103Y112_SLICE_X163Y112_D_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A5Q;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_AMUX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_AO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_AO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_AQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_A_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_BMUX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_BO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_BO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_BQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_B_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_CLK;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_CO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_CO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_CQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_C_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_DO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_DO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_DQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_D_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X162Y113_SR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_AMUX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_AO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_AQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_AX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_A_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_BO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_BO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_BX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_B_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_CLK;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_CO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_CO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_CQ;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_CX;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_C_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D1;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D2;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D3;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D4;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_DO5;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_DO6;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D_CY;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_D_XOR;
  wire [0:0] CLBLM_R_X103Y113_SLICE_X163Y113_SR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_A;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_A1;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_A2;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_A3;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_A4;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_A5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_A6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_AO5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_AO6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_AQ;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_A_CY;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_A_XOR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_B;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_B1;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_B2;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_B3;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_B4;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_B5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_B6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_BO5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_BO6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_BQ;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_B_CY;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_B_XOR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_C;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_C1;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_C2;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_C3;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_C4;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_C5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_C6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_CLK;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_CO5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_CO6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_CQ;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_C_CY;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_C_XOR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_D;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_D1;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_D2;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_D3;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_D4;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_D5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_D6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_DO5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_DO6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_D_CY;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_D_XOR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X162Y114_SR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_A;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_A1;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_A2;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_A3;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_A4;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_A5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_A6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_AO5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_AO6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_AQ;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_A_CY;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_A_XOR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_B;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_B1;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_B2;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_B3;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_B4;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_B5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_B6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_BO5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_BO6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_B_CY;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_B_XOR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_C;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_C1;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_C2;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_C3;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_C4;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_C5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_C6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_CLK;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_CO5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_CO6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_C_CY;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_C_XOR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_D;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_D1;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_D2;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_D3;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_D4;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_D5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_D6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_DO5;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_DO6;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_D_CY;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_D_XOR;
  wire [0:0] CLBLM_R_X103Y114_SLICE_X163Y114_SR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_AMUX;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_AO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_AO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_AQ;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_A_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_BO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_BO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_BQ;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_B_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_CLK;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_CO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_CO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_CQ;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_C_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_DO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_DO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_D_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X162Y115_SR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_AO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_AO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_AQ;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_A_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_BO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_BO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_BQ;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_B_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_CLK;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_CO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_CO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_CQ;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_C_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D1;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D2;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D3;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D4;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_DO5;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_DO6;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_DQ;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D_CY;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_D_XOR;
  wire [0:0] CLBLM_R_X103Y115_SLICE_X163Y115_SR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A5Q;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_AMUX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_AO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_AO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_AQ;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_AX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_A_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B5Q;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_BMUX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_BO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_BO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_BQ;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_BX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_B_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_CLK;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_CO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_CO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_CQ;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_C_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_DMUX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_DO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_D_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X162Y116_SR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A5Q;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_AMUX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_AO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_AO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_AQ;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_A_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B5Q;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_BMUX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_BO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_BO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_BQ;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_BX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_B_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_CLK;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_CMUX;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_CO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_CO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_C_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D1;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D2;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D3;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D4;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_DO5;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_DO6;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_DQ;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D_CY;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_D_XOR;
  wire [0:0] CLBLM_R_X103Y116_SLICE_X163Y116_SR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_AO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_AO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_AQ;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_A_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_BO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_BO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_B_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_CLK;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_CO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_CO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_C_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_DO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_DO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_D_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X162Y117_SR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_AO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_AO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_AQ;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_A_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_BO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_BO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_BQ;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_B_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_CLK;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_CO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_CO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_CQ;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_C_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D1;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D2;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D3;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D4;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_DO5;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_DO6;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D_CY;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_D_XOR;
  wire [0:0] CLBLM_R_X103Y117_SLICE_X163Y117_SR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A1;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A2;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A3;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A4;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_AMUX;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_AO5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_AO6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_AQ;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A_CY;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_A_XOR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B1;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B2;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B3;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B4;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B5Q;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_BMUX;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_BO5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_BO6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_BQ;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_BX;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B_CY;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_B_XOR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_C;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_C1;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_C2;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_C3;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_C4;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_C5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_C6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_CLK;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_CMUX;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_CO5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_CO6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_C_CY;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_C_XOR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_D;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_D1;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_D2;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_D3;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_D4;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_D5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_D6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_DO5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_DO6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_D_CY;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_D_XOR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X162Y118_SR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_A;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_A1;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_A2;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_A3;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_A4;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_A5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_A6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_AO5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_AO6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_AQ;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_AX;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_A_CY;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_A_XOR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_B;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_B1;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_B2;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_B3;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_B4;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_B5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_B6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_BO5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_BO6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_BQ;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_BX;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_B_CY;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_B_XOR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_C;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_C1;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_C2;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_C3;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_C4;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_C5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_C6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_CLK;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_CO5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_CO6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_C_CY;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_C_XOR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_D;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_D1;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_D2;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_D3;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_D4;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_D5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_D6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_DO5;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_DO6;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_D_CY;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_D_XOR;
  wire [0:0] CLBLM_R_X103Y118_SLICE_X163Y118_SR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_AO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_AO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_A_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_BO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_BO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_BQ;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_B_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_CLK;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_CO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_CO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_C_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_DMUX;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_DO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_DO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_D_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X162Y119_SR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_AO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_AO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_A_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_BO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_BO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_B_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_CO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_CO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_C_XOR;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D1;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D2;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D3;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D4;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_DO5;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_DO6;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D_CY;
  wire [0:0] CLBLM_R_X103Y119_SLICE_X163Y119_D_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_A_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_BO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_B_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_CO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_CO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_C_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_DO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X162Y122_D_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_AQ;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_A_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_B_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CLK;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_C_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D1;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D2;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D3;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D4;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_DO5;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D_CY;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_D_XOR;
  wire [0:0] CLBLM_R_X103Y122_SLICE_X163Y122_SR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_O;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_O;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_O;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_O;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_O;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_O;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_O;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_O;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_O;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_O;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_O;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_O;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_O;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_O;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_O;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_O;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_O;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1;
  wire [0:0] RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y115_TQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_D1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_OQ;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_T1;
  wire [0:0] RIOI3_X105Y115_OLOGIC_X1Y116_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y117_TQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_D1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_OQ;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_T1;
  wire [0:0] RIOI3_X105Y117_OLOGIC_X1Y118_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y121_TQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_D1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_OQ;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_T1;
  wire [0:0] RIOI3_X105Y121_OLOGIC_X1Y122_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y123_TQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_D1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_OQ;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_T1;
  wire [0:0] RIOI3_X105Y123_OLOGIC_X1Y124_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y125_TQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_D1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_OQ;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_T1;
  wire [0:0] RIOI3_X105Y125_OLOGIC_X1Y126_TQ;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X105Y127_OLOGIC_X1Y127_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y129_TQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_D1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_OQ;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_T1;
  wire [0:0] RIOI3_X105Y129_OLOGIC_X1Y130_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y133_TQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_D1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_OQ;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_T1;
  wire [0:0] RIOI3_X105Y133_OLOGIC_X1Y134_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y135_TQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_D1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_OQ;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_T1;
  wire [0:0] RIOI3_X105Y135_OLOGIC_X1Y136_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y139_TQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_D1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_OQ;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_T1;
  wire [0:0] RIOI3_X105Y139_OLOGIC_X1Y140_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y141_TQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_D1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_OQ;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_T1;
  wire [0:0] RIOI3_X105Y141_OLOGIC_X1Y142_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y145_TQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_D1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_OQ;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_T1;
  wire [0:0] RIOI3_X105Y145_OLOGIC_X1Y146_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y147_TQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_D1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_OQ;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_T1;
  wire [0:0] RIOI3_X105Y147_OLOGIC_X1Y148_TQ;


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y107_SLICE_X160Y107_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y107_SLICE_X160Y107_AO5),
.Q(CLBLL_L_X102Y107_SLICE_X160Y107_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y107_SLICE_X160Y107_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y107_SLICE_X160Y107_AO6),
.Q(CLBLL_L_X102Y107_SLICE_X160Y107_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y107_SLICE_X160Y107_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y107_SLICE_X160Y107_BO6),
.Q(CLBLL_L_X102Y107_SLICE_X160Y107_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y107_SLICE_X160Y107_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y107_SLICE_X160Y107_CO6),
.Q(CLBLL_L_X102Y107_SLICE_X160Y107_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y107_SLICE_X160Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y107_SLICE_X160Y107_DO5),
.O6(CLBLL_L_X102Y107_SLICE_X160Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffc0003fff)
  ) CLBLL_L_X102Y107_SLICE_X160Y107_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y107_SLICE_X160Y107_AQ),
.I2(CLBLL_L_X102Y107_SLICE_X160Y107_BQ),
.I3(CLBLL_L_X102Y107_SLICE_X160Y107_A5Q),
.I4(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I5(CLBLM_R_X103Y119_SLICE_X162Y119_CO6),
.O5(CLBLL_L_X102Y107_SLICE_X160Y107_CO5),
.O6(CLBLL_L_X102Y107_SLICE_X160Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8808888800800000)
  ) CLBLL_L_X102Y107_SLICE_X160Y107_BLUT (
.I0(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLL_L_X102Y107_SLICE_X160Y107_AQ),
.I3(CLBLM_R_X103Y119_SLICE_X162Y119_CO6),
.I4(CLBLL_L_X102Y107_SLICE_X160Y107_A5Q),
.I5(CLBLL_L_X102Y107_SLICE_X160Y107_BQ),
.O5(CLBLL_L_X102Y107_SLICE_X160Y107_BO5),
.O6(CLBLL_L_X102Y107_SLICE_X160Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8008800888080080)
  ) CLBLL_L_X102Y107_SLICE_X160Y107_ALUT (
.I0(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLL_L_X102Y107_SLICE_X160Y107_AQ),
.I3(CLBLM_R_X103Y119_SLICE_X162Y119_CO6),
.I4(CLBLL_L_X102Y107_SLICE_X160Y107_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y107_SLICE_X160Y107_AO5),
.O6(CLBLL_L_X102Y107_SLICE_X160Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y107_SLICE_X161Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y107_SLICE_X161Y107_DO5),
.O6(CLBLL_L_X102Y107_SLICE_X161Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y107_SLICE_X161Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y107_SLICE_X161Y107_CO5),
.O6(CLBLL_L_X102Y107_SLICE_X161Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y107_SLICE_X161Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y107_SLICE_X161Y107_BO5),
.O6(CLBLL_L_X102Y107_SLICE_X161Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y107_SLICE_X161Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y107_SLICE_X161Y107_AO5),
.O6(CLBLL_L_X102Y107_SLICE_X161Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y108_SLICE_X160Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y108_SLICE_X160Y108_DO5),
.O6(CLBLL_L_X102Y108_SLICE_X160Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y108_SLICE_X160Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y108_SLICE_X160Y108_CO5),
.O6(CLBLL_L_X102Y108_SLICE_X160Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y108_SLICE_X160Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y108_SLICE_X160Y108_BO5),
.O6(CLBLL_L_X102Y108_SLICE_X160Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y108_SLICE_X160Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y108_SLICE_X160Y108_AO5),
.O6(CLBLL_L_X102Y108_SLICE_X160Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y108_SLICE_X161Y108_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y108_SLICE_X161Y108_BO5),
.Q(CLBLL_L_X102Y108_SLICE_X161Y108_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y108_SLICE_X161Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y108_SLICE_X161Y108_AO6),
.Q(CLBLL_L_X102Y108_SLICE_X161Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y108_SLICE_X161Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y108_SLICE_X161Y108_BO6),
.Q(CLBLL_L_X102Y108_SLICE_X161Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y108_SLICE_X161Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y108_SLICE_X161Y108_DO5),
.O6(CLBLL_L_X102Y108_SLICE_X161Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000100)
  ) CLBLL_L_X102Y108_SLICE_X161Y108_CLUT (
.I0(CLBLM_R_X103Y109_SLICE_X163Y109_CQ),
.I1(CLBLL_L_X102Y109_SLICE_X161Y109_AO5),
.I2(CLBLL_L_X102Y108_SLICE_X161Y108_BQ),
.I3(CLBLM_R_X103Y109_SLICE_X162Y109_CQ),
.I4(CLBLL_L_X102Y109_SLICE_X161Y109_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y108_SLICE_X161Y108_CO5),
.O6(CLBLL_L_X102Y108_SLICE_X161Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c050505050)
  ) CLBLL_L_X102Y108_SLICE_X161Y108_BLUT (
.I0(CLBLM_R_X103Y109_SLICE_X162Y109_CQ),
.I1(CLBLL_L_X102Y110_SLICE_X161Y110_B5Q),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y108_SLICE_X161Y108_BO5),
.O6(CLBLL_L_X102Y108_SLICE_X161Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0d0d0c0c0c0c0)
  ) CLBLL_L_X102Y108_SLICE_X161Y108_ALUT (
.I0(CLBLL_L_X102Y109_SLICE_X161Y109_DO6),
.I1(CLBLL_L_X102Y109_SLICE_X161Y109_CO5),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(CLBLM_R_X103Y109_SLICE_X162Y109_DO6),
.I5(CLBLL_L_X102Y108_SLICE_X161Y108_CO6),
.O5(CLBLL_L_X102Y108_SLICE_X161Y108_AO5),
.O6(CLBLL_L_X102Y108_SLICE_X161Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X160Y109_AO5),
.Q(CLBLL_L_X102Y109_SLICE_X160Y109_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X160Y109_BO5),
.Q(CLBLL_L_X102Y109_SLICE_X160Y109_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X160Y109_CO5),
.Q(CLBLL_L_X102Y109_SLICE_X160Y109_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X160Y109_AO6),
.Q(CLBLL_L_X102Y109_SLICE_X160Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X160Y109_BO6),
.Q(CLBLL_L_X102Y109_SLICE_X160Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X160Y109_CO6),
.Q(CLBLL_L_X102Y109_SLICE_X160Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y109_SLICE_X160Y109_DO5),
.O6(CLBLL_L_X102Y109_SLICE_X160Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff003333)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y109_SLICE_X160Y109_AQ),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLL_L_X102Y109_SLICE_X161Y109_CQ),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X102Y109_SLICE_X160Y109_CO5),
.O6(CLBLL_L_X102Y109_SLICE_X160Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0000050505050)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_BLUT (
.I0(CLBLM_R_X103Y112_SLICE_X162Y112_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(CLBLL_L_X102Y108_SLICE_X161Y108_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y109_SLICE_X160Y109_BO5),
.O6(CLBLL_L_X102Y109_SLICE_X160Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff55ffe4ffe4)
  ) CLBLL_L_X102Y109_SLICE_X160Y109_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLL_L_X102Y110_SLICE_X160Y110_D5Q),
.I2(CLBLL_L_X102Y109_SLICE_X161Y109_B5Q),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I4(CLBLL_L_X102Y109_SLICE_X161Y109_CQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y109_SLICE_X160Y109_AO5),
.O6(CLBLL_L_X102Y109_SLICE_X160Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X161Y109_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X161Y109_BO5),
.Q(CLBLL_L_X102Y109_SLICE_X161Y109_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X161Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X161Y109_AO6),
.Q(CLBLL_L_X102Y109_SLICE_X161Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X161Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X161Y109_BO6),
.Q(CLBLL_L_X102Y109_SLICE_X161Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X161Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X161Y109_CO6),
.Q(CLBLL_L_X102Y109_SLICE_X161Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y109_SLICE_X161Y109_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y109_SLICE_X160Y109_C5Q),
.Q(CLBLL_L_X102Y109_SLICE_X161Y109_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff3f)
  ) CLBLL_L_X102Y109_SLICE_X161Y109_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y108_SLICE_X162Y108_BQ),
.I2(CLBLM_R_X103Y112_SLICE_X162Y112_AQ),
.I3(CLBLL_L_X102Y109_SLICE_X160Y109_CQ),
.I4(CLBLM_R_X103Y109_SLICE_X163Y109_CO6),
.I5(CLBLL_L_X102Y109_SLICE_X160Y109_BQ),
.O5(CLBLL_L_X102Y109_SLICE_X161Y109_DO5),
.O6(CLBLL_L_X102Y109_SLICE_X161Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000069966996)
  ) CLBLL_L_X102Y109_SLICE_X161Y109_CLUT (
.I0(CLBLL_L_X102Y108_SLICE_X161Y108_AQ),
.I1(CLBLL_L_X102Y109_SLICE_X161Y109_AQ),
.I2(CLBLM_R_X103Y109_SLICE_X162Y109_AQ),
.I3(CLBLL_L_X102Y110_SLICE_X161Y110_BQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X102Y109_SLICE_X161Y109_CO5),
.O6(CLBLL_L_X102Y109_SLICE_X161Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLL_L_X102Y109_SLICE_X161Y109_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y109_SLICE_X160Y109_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLL_L_X102Y108_SLICE_X161Y108_AQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y109_SLICE_X161Y109_BO5),
.O6(CLBLL_L_X102Y109_SLICE_X161Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fffbfffb)
  ) CLBLL_L_X102Y109_SLICE_X161Y109_ALUT (
.I0(CLBLL_L_X102Y110_SLICE_X161Y110_BQ),
.I1(CLBLL_L_X102Y109_SLICE_X160Y109_B5Q),
.I2(CLBLL_L_X102Y108_SLICE_X161Y108_AQ),
.I3(CLBLL_L_X102Y109_SLICE_X161Y109_CQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X102Y109_SLICE_X161Y109_AO5),
.O6(CLBLL_L_X102Y109_SLICE_X161Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_AO5),
.Q(CLBLL_L_X102Y110_SLICE_X160Y110_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_BO5),
.Q(CLBLL_L_X102Y110_SLICE_X160Y110_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_CO5),
.Q(CLBLL_L_X102Y110_SLICE_X160Y110_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_DO5),
.Q(CLBLL_L_X102Y110_SLICE_X160Y110_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_AO6),
.Q(CLBLL_L_X102Y110_SLICE_X160Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_BO6),
.Q(CLBLL_L_X102Y110_SLICE_X160Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_CO6),
.Q(CLBLL_L_X102Y110_SLICE_X160Y110_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_DO6),
.Q(CLBLL_L_X102Y110_SLICE_X160Y110_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa000000aaaa)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X103Y109_SLICE_X162Y109_A5Q),
.I4(CLBLL_L_X102Y109_SLICE_X160Y109_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y110_SLICE_X160Y110_DO5),
.O6(CLBLL_L_X102Y110_SLICE_X160Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dd110000cf03)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_CLUT (
.I0(CLBLL_L_X102Y110_SLICE_X160Y110_C5Q),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLL_L_X102Y110_SLICE_X160Y110_BQ),
.I3(CLBLM_R_X103Y109_SLICE_X162Y109_A5Q),
.I4(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y110_SLICE_X160Y110_CO5),
.O6(CLBLL_L_X102Y110_SLICE_X160Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000aaaa3333)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_BLUT (
.I0(CLBLL_L_X102Y109_SLICE_X161Y109_B5Q),
.I1(CLBLL_L_X102Y109_SLICE_X160Y109_A5Q),
.I2(CLBLL_L_X102Y109_SLICE_X160Y109_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X102Y110_SLICE_X160Y110_BO5),
.O6(CLBLL_L_X102Y110_SLICE_X160Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0333350500055)
  ) CLBLL_L_X102Y110_SLICE_X160Y110_ALUT (
.I0(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I1(CLBLL_L_X102Y110_SLICE_X160Y110_A5Q),
.I2(CLBLL_L_X102Y109_SLICE_X160Y109_BQ),
.I3(CLBLM_R_X103Y110_SLICE_X162Y110_AQ),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X102Y110_SLICE_X160Y110_AO5),
.O6(CLBLL_L_X102Y110_SLICE_X160Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X161Y110_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X161Y110_AO5),
.Q(CLBLL_L_X102Y110_SLICE_X161Y110_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X161Y110_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X161Y110_BO5),
.Q(CLBLL_L_X102Y110_SLICE_X161Y110_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X161Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X161Y110_AO6),
.Q(CLBLL_L_X102Y110_SLICE_X161Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X161Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X161Y110_BO6),
.Q(CLBLL_L_X102Y110_SLICE_X161Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y110_SLICE_X161Y110_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y111_SLICE_X161Y111_DQ),
.Q(CLBLL_L_X102Y110_SLICE_X161Y110_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y110_SLICE_X161Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y110_SLICE_X161Y110_DO5),
.O6(CLBLL_L_X102Y110_SLICE_X161Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y110_SLICE_X161Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y110_SLICE_X161Y110_CO5),
.O6(CLBLL_L_X102Y110_SLICE_X161Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X102Y110_SLICE_X161Y110_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLL_L_X102Y109_SLICE_X161Y109_BQ),
.I2(CLBLM_R_X103Y109_SLICE_X162Y109_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y110_SLICE_X161Y110_BO5),
.O6(CLBLL_L_X102Y110_SLICE_X161Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3030300f50005)
  ) CLBLL_L_X102Y110_SLICE_X161Y110_ALUT (
.I0(CLBLL_L_X102Y110_SLICE_X160Y110_DQ),
.I1(CLBLL_L_X102Y110_SLICE_X161Y110_A5Q),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I4(CLBLM_R_X103Y109_SLICE_X163Y109_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y110_SLICE_X161Y110_AO5),
.O6(CLBLL_L_X102Y110_SLICE_X161Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_DQ),
.Q(CLBLL_L_X102Y111_SLICE_X160Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_A5Q),
.Q(CLBLL_L_X102Y111_SLICE_X160Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X161Y110_CQ),
.Q(CLBLL_L_X102Y111_SLICE_X160Y111_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_AO5),
.Q(CLBLL_L_X102Y111_SLICE_X160Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_BO5),
.Q(CLBLL_L_X102Y111_SLICE_X160Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_CO5),
.Q(CLBLL_L_X102Y111_SLICE_X160Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_CQ),
.Q(CLBLL_L_X102Y111_SLICE_X160Y111_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0ff0e00f0e)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_DLUT (
.I0(CLBLL_L_X102Y111_SLICE_X160Y111_AO6),
.I1(CLBLL_L_X102Y112_SLICE_X160Y112_CO6),
.I2(CLBLL_L_X102Y112_SLICE_X160Y112_B5Q),
.I3(CLBLL_L_X102Y111_SLICE_X160Y111_CO6),
.I4(CLBLL_L_X102Y112_SLICE_X160Y112_CQ),
.I5(CLBLL_L_X102Y111_SLICE_X160Y111_BO6),
.O5(CLBLL_L_X102Y111_SLICE_X160Y111_DO5),
.O6(CLBLL_L_X102Y111_SLICE_X160Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffcffff0000)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y112_SLICE_X160Y112_A5Q),
.I2(CLBLL_L_X102Y112_SLICE_X160Y112_B5Q),
.I3(CLBLL_L_X102Y110_SLICE_X161Y110_CQ),
.I4(CLBLL_L_X102Y111_SLICE_X160Y111_BQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y111_SLICE_X160Y111_CO5),
.O6(CLBLL_L_X102Y111_SLICE_X160Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefeff00ff00)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_BLUT (
.I0(CLBLL_L_X102Y112_SLICE_X161Y112_B5Q),
.I1(CLBLL_L_X102Y111_SLICE_X160Y111_A5Q),
.I2(CLBLL_L_X102Y111_SLICE_X160Y111_DQ),
.I3(CLBLL_L_X102Y112_SLICE_X160Y112_A5Q),
.I4(CLBLL_L_X102Y111_SLICE_X160Y111_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X102Y111_SLICE_X160Y111_BO5),
.O6(CLBLL_L_X102Y111_SLICE_X160Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefeff00ff00)
  ) CLBLL_L_X102Y111_SLICE_X160Y111_ALUT (
.I0(CLBLL_L_X102Y112_SLICE_X160Y112_CQ),
.I1(CLBLL_L_X102Y111_SLICE_X160Y111_BQ),
.I2(CLBLL_L_X102Y111_SLICE_X161Y111_DQ),
.I3(CLBLL_L_X102Y110_SLICE_X160Y110_B5Q),
.I4(CLBLL_L_X102Y112_SLICE_X161Y112_AQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y111_SLICE_X160Y111_AO5),
.O6(CLBLL_L_X102Y111_SLICE_X160Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_CQ),
.Q(CLBLL_L_X102Y111_SLICE_X161Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y111_SLICE_X162Y111_BQ),
.Q(CLBLL_L_X102Y111_SLICE_X161Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X161Y110_AQ),
.Q(CLBLL_L_X102Y111_SLICE_X161Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y112_SLICE_X161Y112_B5Q),
.Q(CLBLL_L_X102Y111_SLICE_X161Y111_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffc3ffc3ffff)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y111_SLICE_X163Y111_DQ),
.I2(CLBLL_L_X102Y111_SLICE_X160Y111_B5Q),
.I3(CLBLL_L_X102Y111_SLICE_X161Y111_CO6),
.I4(CLBLL_L_X102Y109_SLICE_X161Y109_DQ),
.I5(CLBLL_L_X102Y111_SLICE_X161Y111_DQ),
.O5(CLBLL_L_X102Y111_SLICE_X161Y111_DO5),
.O6(CLBLL_L_X102Y111_SLICE_X161Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hebffd7ffffebffd7)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_CLUT (
.I0(CLBLL_L_X102Y111_SLICE_X160Y111_AQ),
.I1(CLBLL_L_X102Y111_SLICE_X160Y111_A5Q),
.I2(CLBLM_R_X103Y111_SLICE_X163Y111_CQ),
.I3(CLBLL_L_X102Y112_SLICE_X161Y112_AQ),
.I4(CLBLL_L_X102Y112_SLICE_X161Y112_B5Q),
.I5(CLBLM_R_X103Y111_SLICE_X163Y111_AQ),
.O5(CLBLL_L_X102Y111_SLICE_X161Y111_CO5),
.O6(CLBLL_L_X102Y111_SLICE_X161Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00eeee0000e0e000)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_BLUT (
.I0(CLBLL_L_X102Y111_SLICE_X161Y111_AQ),
.I1(CLBLL_L_X102Y112_SLICE_X160Y112_A5Q),
.I2(CLBLL_L_X102Y111_SLICE_X161Y111_CQ),
.I3(CLBLL_L_X102Y111_SLICE_X160Y111_DQ),
.I4(CLBLM_R_X103Y111_SLICE_X163Y111_BQ),
.I5(CLBLL_L_X102Y111_SLICE_X160Y111_CQ),
.O5(CLBLL_L_X102Y111_SLICE_X161Y111_BO5),
.O6(CLBLL_L_X102Y111_SLICE_X161Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefbeebbfcf3cc33)
  ) CLBLL_L_X102Y111_SLICE_X161Y111_ALUT (
.I0(CLBLL_L_X102Y111_SLICE_X161Y111_AQ),
.I1(CLBLL_L_X102Y111_SLICE_X161Y111_BQ),
.I2(CLBLL_L_X102Y111_SLICE_X161Y111_CQ),
.I3(CLBLL_L_X102Y111_SLICE_X160Y111_BQ),
.I4(CLBLL_L_X102Y111_SLICE_X160Y111_CQ),
.I5(CLBLL_L_X102Y112_SLICE_X160Y112_A5Q),
.O5(CLBLL_L_X102Y111_SLICE_X161Y111_AO5),
.O6(CLBLL_L_X102Y111_SLICE_X161Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y112_SLICE_X161Y112_AQ),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y112_SLICE_X160Y112_CQ),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_C5Q),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y112_SLICE_X160Y112_AO6),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y112_SLICE_X160Y112_BO6),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y112_SLICE_X160Y112_CO5),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y112_SLICE_X160Y112_C5Q),
.Q(CLBLL_L_X102Y112_SLICE_X160Y112_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y112_SLICE_X160Y112_DO5),
.O6(CLBLL_L_X102Y112_SLICE_X160Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffef0f0f0f0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_CLUT (
.I0(CLBLL_L_X102Y112_SLICE_X160Y112_C5Q),
.I1(CLBLL_L_X102Y111_SLICE_X160Y111_CQ),
.I2(CLBLL_L_X102Y112_SLICE_X160Y112_DQ),
.I3(CLBLL_L_X102Y111_SLICE_X160Y111_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y112_SLICE_X160Y112_CO5),
.O6(CLBLL_L_X102Y112_SLICE_X160Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a8888888)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLL_L_X102Y112_SLICE_X160Y112_BQ),
.I2(CLBLL_L_X102Y112_SLICE_X160Y112_AQ),
.I3(CLBLL_L_X102Y112_SLICE_X161Y112_BQ),
.I4(CLBLL_L_X102Y113_SLICE_X161Y113_AQ),
.I5(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.O5(CLBLL_L_X102Y112_SLICE_X160Y112_BO5),
.O6(CLBLL_L_X102Y112_SLICE_X160Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000008aa0a0a0)
  ) CLBLL_L_X102Y112_SLICE_X160Y112_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLL_L_X102Y112_SLICE_X160Y112_BQ),
.I2(CLBLL_L_X102Y112_SLICE_X160Y112_AQ),
.I3(CLBLL_L_X102Y112_SLICE_X161Y112_BQ),
.I4(CLBLL_L_X102Y113_SLICE_X161Y113_AQ),
.I5(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.O5(CLBLL_L_X102Y112_SLICE_X160Y112_AO5),
.O6(CLBLL_L_X102Y112_SLICE_X160Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y110_SLICE_X160Y110_AQ),
.Q(CLBLL_L_X102Y112_SLICE_X161Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y111_SLICE_X160Y111_B5Q),
.Q(CLBLL_L_X102Y112_SLICE_X161Y112_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y112_SLICE_X161Y112_AO6),
.Q(CLBLL_L_X102Y112_SLICE_X161Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y112_SLICE_X161Y112_BO6),
.Q(CLBLL_L_X102Y112_SLICE_X161Y112_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3fffffffffffff)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y113_SLICE_X161Y113_AQ),
.I2(CLBLL_L_X102Y112_SLICE_X161Y112_BQ),
.I3(1'b1),
.I4(CLBLL_L_X102Y112_SLICE_X160Y112_AQ),
.I5(CLBLL_L_X102Y112_SLICE_X160Y112_BQ),
.O5(CLBLL_L_X102Y112_SLICE_X161Y112_DO5),
.O6(CLBLL_L_X102Y112_SLICE_X161Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0110ffff0000)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_CLUT (
.I0(CLBLL_L_X102Y111_SLICE_X161Y111_AO6),
.I1(CLBLL_L_X102Y111_SLICE_X161Y111_DO6),
.I2(CLBLL_L_X102Y111_SLICE_X160Y111_DO6),
.I3(CLBLL_L_X102Y112_SLICE_X161Y112_A5Q),
.I4(CLBLL_L_X102Y112_SLICE_X161Y112_DO6),
.I5(CLBLL_L_X102Y111_SLICE_X161Y111_BO6),
.O5(CLBLL_L_X102Y112_SLICE_X161Y112_CO5),
.O6(CLBLL_L_X102Y112_SLICE_X161Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a2222222)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLL_L_X102Y112_SLICE_X161Y112_BQ),
.I2(CLBLL_L_X102Y113_SLICE_X161Y113_AQ),
.I3(CLBLL_L_X102Y112_SLICE_X160Y112_BQ),
.I4(CLBLL_L_X102Y112_SLICE_X160Y112_AQ),
.I5(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.O5(CLBLL_L_X102Y112_SLICE_X161Y112_BO5),
.O6(CLBLL_L_X102Y112_SLICE_X161Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff40000000)
  ) CLBLL_L_X102Y112_SLICE_X161Y112_ALUT (
.I0(CLBLL_L_X102Y111_SLICE_X160Y111_DO6),
.I1(CLBLL_L_X102Y112_SLICE_X161Y112_BQ),
.I2(CLBLL_L_X102Y113_SLICE_X161Y113_AQ),
.I3(CLBLL_L_X102Y112_SLICE_X160Y112_BQ),
.I4(CLBLL_L_X102Y112_SLICE_X160Y112_AQ),
.I5(CLBLL_L_X102Y112_SLICE_X161Y112_A5Q),
.O5(CLBLL_L_X102Y112_SLICE_X161Y112_AO5),
.O6(CLBLL_L_X102Y112_SLICE_X161Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X160Y113_DO5),
.O6(CLBLL_L_X102Y113_SLICE_X160Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X160Y113_CO5),
.O6(CLBLL_L_X102Y113_SLICE_X160Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X160Y113_BO5),
.O6(CLBLL_L_X102Y113_SLICE_X160Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X160Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X160Y113_AO5),
.O6(CLBLL_L_X102Y113_SLICE_X160Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y113_SLICE_X161Y113_AO6),
.Q(CLBLL_L_X102Y113_SLICE_X161Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X161Y113_DO5),
.O6(CLBLL_L_X102Y113_SLICE_X161Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X161Y113_CO5),
.O6(CLBLL_L_X102Y113_SLICE_X161Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y113_SLICE_X161Y113_BO5),
.O6(CLBLL_L_X102Y113_SLICE_X161Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000c8484848)
  ) CLBLL_L_X102Y113_SLICE_X161Y113_ALUT (
.I0(CLBLL_L_X102Y113_SLICE_X161Y113_AQ),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLL_L_X102Y112_SLICE_X161Y112_BQ),
.I3(CLBLL_L_X102Y112_SLICE_X160Y112_BQ),
.I4(CLBLL_L_X102Y112_SLICE_X160Y112_AQ),
.I5(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.O5(CLBLL_L_X102Y113_SLICE_X161Y113_AO5),
.O6(CLBLL_L_X102Y113_SLICE_X161Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X160Y114_DO5),
.O6(CLBLL_L_X102Y114_SLICE_X160Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X160Y114_CO5),
.O6(CLBLL_L_X102Y114_SLICE_X160Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X160Y114_BO5),
.O6(CLBLL_L_X102Y114_SLICE_X160Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X160Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X160Y114_AO5),
.O6(CLBLL_L_X102Y114_SLICE_X160Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y114_SLICE_X161Y114_AO6),
.Q(CLBLL_L_X102Y114_SLICE_X161Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X161Y114_DO5),
.O6(CLBLL_L_X102Y114_SLICE_X161Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X161Y114_CO5),
.O6(CLBLL_L_X102Y114_SLICE_X161Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y114_SLICE_X161Y114_BO5),
.O6(CLBLL_L_X102Y114_SLICE_X161Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0cc00ccf0f00000)
  ) CLBLL_L_X102Y114_SLICE_X161Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y114_SLICE_X162Y114_CQ),
.I2(CLBLL_L_X102Y114_SLICE_X161Y114_AQ),
.I3(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.O5(CLBLL_L_X102Y114_SLICE_X161Y114_AO5),
.O6(CLBLL_L_X102Y114_SLICE_X161Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y115_SLICE_X160Y115_AO6),
.Q(CLBLL_L_X102Y115_SLICE_X160Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y115_SLICE_X160Y115_DO5),
.O6(CLBLL_L_X102Y115_SLICE_X160Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y115_SLICE_X160Y115_CO5),
.O6(CLBLL_L_X102Y115_SLICE_X160Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X102Y115_SLICE_X160Y115_BO5),
.O6(CLBLL_L_X102Y115_SLICE_X160Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0eac0eac040c040)
  ) CLBLL_L_X102Y115_SLICE_X160Y115_ALUT (
.I0(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLL_L_X102Y115_SLICE_X160Y115_AQ),
.I3(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I4(1'b1),
.I5(CLBLL_L_X102Y115_SLICE_X161Y115_CQ),
.O5(CLBLL_L_X102Y115_SLICE_X160Y115_AO5),
.O6(CLBLL_L_X102Y115_SLICE_X160Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.Q(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y115_SLICE_X161Y115_AO6),
.Q(CLBLL_L_X102Y115_SLICE_X161Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y115_SLICE_X161Y115_BO6),
.Q(CLBLL_L_X102Y115_SLICE_X161Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLL_L_X102Y115_SLICE_X161Y115_CO6),
.Q(CLBLL_L_X102Y115_SLICE_X161Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffee)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_DLUT (
.I0(CLBLL_L_X102Y115_SLICE_X160Y115_AQ),
.I1(CLBLL_L_X102Y115_SLICE_X161Y115_CQ),
.I2(1'b1),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_BQ),
.I4(CLBLL_L_X102Y115_SLICE_X161Y115_AQ),
.I5(CLBLM_R_X103Y116_SLICE_X162Y116_BQ),
.O5(CLBLL_L_X102Y115_SLICE_X161Y115_DO5),
.O6(CLBLL_L_X102Y115_SLICE_X161Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc50dc508c008c00)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_CLUT (
.I0(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I1(CLBLL_L_X102Y115_SLICE_X161Y115_CQ),
.I2(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(CLBLM_R_X103Y115_SLICE_X162Y115_CQ),
.O5(CLBLL_L_X102Y115_SLICE_X161Y115_CO5),
.O6(CLBLL_L_X102Y115_SLICE_X161Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hce0ac400ce0ac400)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_BLUT (
.I0(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I1(CLBLL_L_X102Y115_SLICE_X161Y115_BQ),
.I2(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLL_L_X102Y115_SLICE_X160Y115_AQ),
.I5(1'b1),
.O5(CLBLL_L_X102Y115_SLICE_X161Y115_BO5),
.O6(CLBLL_L_X102Y115_SLICE_X161Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd08fd0808080808)
  ) CLBLL_L_X102Y115_SLICE_X161Y115_ALUT (
.I0(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I1(CLBLL_L_X102Y115_SLICE_X161Y115_BQ),
.I2(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(CLBLL_L_X102Y115_SLICE_X161Y115_AQ),
.O5(CLBLL_L_X102Y115_SLICE_X161Y115_AO5),
.O6(CLBLL_L_X102Y115_SLICE_X161Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y108_SLICE_X162Y108_AO5),
.Q(CLBLM_R_X103Y108_SLICE_X162Y108_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y108_SLICE_X162Y108_BO5),
.Q(CLBLM_R_X103Y108_SLICE_X162Y108_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y108_SLICE_X162Y108_AO6),
.Q(CLBLM_R_X103Y108_SLICE_X162Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y108_SLICE_X162Y108_BO6),
.Q(CLBLM_R_X103Y108_SLICE_X162Y108_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_DO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0000000ff0000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(1'b1),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X103Y109_SLICE_X163Y109_AQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_CO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000f0f00000)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(1'b1),
.I4(CLBLM_R_X103Y108_SLICE_X163Y108_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_BO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ff330d010d01)
  ) CLBLM_R_X103Y108_SLICE_X162Y108_ALUT (
.I0(CLBLM_R_X103Y108_SLICE_X162Y108_B5Q),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I3(CLBLM_R_X103Y109_SLICE_X163Y109_CQ),
.I4(CLBLM_R_X103Y108_SLICE_X162Y108_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X162Y108_AO5),
.O6(CLBLM_R_X103Y108_SLICE_X162Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y108_SLICE_X162Y108_CO5),
.Q(CLBLM_R_X103Y108_SLICE_X163Y108_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_DO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_CO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_BO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y108_SLICE_X163Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y108_SLICE_X163Y108_AO5),
.O6(CLBLM_R_X103Y108_SLICE_X163Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y109_SLICE_X162Y109_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y109_SLICE_X162Y109_AO5),
.Q(CLBLM_R_X103Y109_SLICE_X162Y109_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y109_SLICE_X162Y109_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y109_SLICE_X162Y109_BO5),
.Q(CLBLM_R_X103Y109_SLICE_X162Y109_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y109_SLICE_X162Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y109_SLICE_X162Y109_AO6),
.Q(CLBLM_R_X103Y109_SLICE_X162Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y109_SLICE_X162Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y109_SLICE_X162Y109_BO6),
.Q(CLBLM_R_X103Y109_SLICE_X162Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y109_SLICE_X162Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y109_SLICE_X162Y109_CO6),
.Q(CLBLM_R_X103Y109_SLICE_X162Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffee)
  ) CLBLM_R_X103Y109_SLICE_X162Y109_DLUT (
.I0(CLBLM_R_X103Y109_SLICE_X162Y109_CO5),
.I1(CLBLL_L_X102Y110_SLICE_X161Y110_B5Q),
.I2(1'b1),
.I3(CLBLM_R_X103Y109_SLICE_X162Y109_A5Q),
.I4(CLBLM_R_X103Y108_SLICE_X163Y108_AQ),
.I5(CLBLM_R_X103Y109_SLICE_X163Y109_BQ),
.O5(CLBLM_R_X103Y109_SLICE_X162Y109_DO5),
.O6(CLBLM_R_X103Y109_SLICE_X162Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ffffffdd)
  ) CLBLM_R_X103Y109_SLICE_X162Y109_CLUT (
.I0(CLBLM_R_X103Y109_SLICE_X163Y109_AQ),
.I1(CLBLM_R_X103Y109_SLICE_X162Y109_AQ),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLL_L_X102Y109_SLICE_X161Y109_B5Q),
.I4(CLBLM_R_X103Y109_SLICE_X162Y109_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y109_SLICE_X162Y109_CO5),
.O6(CLBLM_R_X103Y109_SLICE_X162Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550000cccc0000)
  ) CLBLM_R_X103Y109_SLICE_X162Y109_BLUT (
.I0(CLBLL_L_X102Y109_SLICE_X160Y109_B5Q),
.I1(CLBLM_R_X103Y109_SLICE_X162Y109_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y109_SLICE_X162Y109_BO5),
.O6(CLBLM_R_X103Y109_SLICE_X162Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0000033330000)
  ) CLBLM_R_X103Y109_SLICE_X162Y109_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y108_SLICE_X162Y108_BQ),
.I2(CLBLL_L_X102Y109_SLICE_X160Y109_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y109_SLICE_X162Y109_AO5),
.O6(CLBLM_R_X103Y109_SLICE_X162Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y109_SLICE_X163Y109_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y109_SLICE_X163Y109_BO5),
.Q(CLBLM_R_X103Y109_SLICE_X163Y109_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y109_SLICE_X163Y109_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y109_SLICE_X163Y109_AO6),
.Q(CLBLM_R_X103Y109_SLICE_X163Y109_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y109_SLICE_X163Y109_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y109_SLICE_X163Y109_BO6),
.Q(CLBLM_R_X103Y109_SLICE_X163Y109_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y109_SLICE_X163Y109_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y109_SLICE_X163Y109_CO5),
.Q(CLBLM_R_X103Y109_SLICE_X163Y109_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y109_SLICE_X163Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y109_SLICE_X163Y109_DO5),
.O6(CLBLM_R_X103Y109_SLICE_X163Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdfdf0f000f00)
  ) CLBLM_R_X103Y109_SLICE_X163Y109_CLUT (
.I0(CLBLL_L_X102Y108_SLICE_X161Y108_B5Q),
.I1(CLBLL_L_X102Y109_SLICE_X161Y109_AQ),
.I2(CLBLM_R_X103Y109_SLICE_X162Y109_BQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X103Y109_SLICE_X163Y109_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y109_SLICE_X163Y109_CO5),
.O6(CLBLM_R_X103Y109_SLICE_X163Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0c0c0c0c0)
  ) CLBLM_R_X103Y109_SLICE_X163Y109_BLUT (
.I0(CLBLM_R_X103Y109_SLICE_X163Y109_CQ),
.I1(CLBLM_R_X103Y109_SLICE_X163Y109_BQ),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y109_SLICE_X163Y109_BO5),
.O6(CLBLM_R_X103Y109_SLICE_X163Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0c000c000)
  ) CLBLM_R_X103Y109_SLICE_X163Y109_ALUT (
.I0(CLBLM_R_X103Y109_SLICE_X163Y109_B5Q),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y109_SLICE_X163Y109_AO5),
.O6(CLBLM_R_X103Y109_SLICE_X163Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_AO5),
.Q(CLBLM_R_X103Y110_SLICE_X162Y110_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_BO5),
.Q(CLBLM_R_X103Y110_SLICE_X162Y110_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_C5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_CO5),
.Q(CLBLM_R_X103Y110_SLICE_X162Y110_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_D5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_DO5),
.Q(CLBLM_R_X103Y110_SLICE_X162Y110_D5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_AO6),
.Q(CLBLM_R_X103Y110_SLICE_X162Y110_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_BO6),
.Q(CLBLM_R_X103Y110_SLICE_X162Y110_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_CO6),
.Q(CLBLM_R_X103Y110_SLICE_X162Y110_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_DO6),
.Q(CLBLM_R_X103Y110_SLICE_X162Y110_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a5f5f001b001b)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_R_X103Y110_SLICE_X162Y110_CQ),
.I2(CLBLL_L_X102Y109_SLICE_X160Y109_B5Q),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I4(CLBLM_R_X103Y110_SLICE_X162Y110_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y110_SLICE_X162Y110_DO5),
.O6(CLBLM_R_X103Y110_SLICE_X162Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000aaaa0000)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_CLUT (
.I0(CLBLM_R_X103Y109_SLICE_X163Y109_CQ),
.I1(1'b1),
.I2(CLBLM_R_X103Y109_SLICE_X163Y109_B5Q),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y110_SLICE_X162Y110_CO5),
.O6(CLBLM_R_X103Y110_SLICE_X162Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbffbbaeaebfbf)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_BLUT (
.I0(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLL_L_X102Y108_SLICE_X161Y108_B5Q),
.I3(CLBLL_L_X102Y110_SLICE_X161Y110_B5Q),
.I4(CLBLM_R_X103Y110_SLICE_X162Y110_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y110_SLICE_X162Y110_BO5),
.O6(CLBLM_R_X103Y110_SLICE_X162Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff000f550f55)
  ) CLBLM_R_X103Y110_SLICE_X162Y110_ALUT (
.I0(CLBLM_R_X103Y110_SLICE_X162Y110_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X102Y108_SLICE_X161Y108_B5Q),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLL_L_X102Y108_SLICE_X161Y108_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y110_SLICE_X162Y110_AO5),
.O6(CLBLM_R_X103Y110_SLICE_X162Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y110_SLICE_X163Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y110_SLICE_X163Y110_DO5),
.O6(CLBLM_R_X103Y110_SLICE_X163Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y110_SLICE_X163Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y110_SLICE_X163Y110_CO5),
.O6(CLBLM_R_X103Y110_SLICE_X163Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y110_SLICE_X163Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y110_SLICE_X163Y110_BO5),
.O6(CLBLM_R_X103Y110_SLICE_X163Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y110_SLICE_X163Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y110_SLICE_X163Y110_AO5),
.O6(CLBLM_R_X103Y110_SLICE_X163Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y111_SLICE_X162Y111_AO5),
.Q(CLBLM_R_X103Y111_SLICE_X162Y111_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y111_SLICE_X162Y111_BO5),
.Q(CLBLM_R_X103Y111_SLICE_X162Y111_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y111_SLICE_X162Y111_AO6),
.Q(CLBLM_R_X103Y111_SLICE_X162Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y111_SLICE_X162Y111_BO6),
.Q(CLBLM_R_X103Y111_SLICE_X162Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X162Y111_DO5),
.O6(CLBLM_R_X103Y111_SLICE_X162Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X162Y111_CO5),
.O6(CLBLM_R_X103Y111_SLICE_X162Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00555533000303)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_BLUT (
.I0(CLBLM_R_X103Y111_SLICE_X162Y111_B5Q),
.I1(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I2(CLBLM_R_X103Y111_SLICE_X162Y111_AQ),
.I3(CLBLM_R_X103Y108_SLICE_X163Y108_AQ),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X162Y111_BO5),
.O6(CLBLM_R_X103Y111_SLICE_X162Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cccc00ff)
  ) CLBLM_R_X103Y111_SLICE_X162Y111_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X102Y110_SLICE_X161Y110_B5Q),
.I2(1'b1),
.I3(CLBLM_R_X103Y110_SLICE_X162Y110_BQ),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X162Y111_AO5),
.O6(CLBLM_R_X103Y111_SLICE_X162Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y111_SLICE_X162Y111_A5Q),
.Q(CLBLM_R_X103Y111_SLICE_X163Y111_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y108_SLICE_X162Y108_AQ),
.Q(CLBLM_R_X103Y111_SLICE_X163Y111_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_DQ),
.Q(CLBLM_R_X103Y111_SLICE_X163Y111_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y110_SLICE_X162Y110_A5Q),
.Q(CLBLM_R_X103Y111_SLICE_X163Y111_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X163Y111_DO5),
.O6(CLBLM_R_X103Y111_SLICE_X163Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X163Y111_CO5),
.O6(CLBLM_R_X103Y111_SLICE_X163Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X163Y111_BO5),
.O6(CLBLM_R_X103Y111_SLICE_X163Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y111_SLICE_X163Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y111_SLICE_X163Y111_AO5),
.O6(CLBLM_R_X103Y111_SLICE_X163Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y112_SLICE_X162Y112_AO5),
.Q(CLBLM_R_X103Y112_SLICE_X162Y112_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y112_SLICE_X162Y112_AO6),
.Q(CLBLM_R_X103Y112_SLICE_X162Y112_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X162Y112_DO5),
.O6(CLBLM_R_X103Y112_SLICE_X162Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X162Y112_CO5),
.O6(CLBLM_R_X103Y112_SLICE_X162Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X162Y112_BO5),
.O6(CLBLM_R_X103Y112_SLICE_X162Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff0022002200)
  ) CLBLM_R_X103Y112_SLICE_X162Y112_ALUT (
.I0(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I1(CLBLM_R_X103Y112_SLICE_X162Y112_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLL_L_X102Y108_SLICE_X161Y108_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X162Y112_AO5),
.O6(CLBLM_R_X103Y112_SLICE_X162Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X163Y112_DO5),
.O6(CLBLM_R_X103Y112_SLICE_X163Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X163Y112_CO5),
.O6(CLBLM_R_X103Y112_SLICE_X163Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X163Y112_BO5),
.O6(CLBLM_R_X103Y112_SLICE_X163Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y112_SLICE_X163Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y112_SLICE_X163Y112_AO5),
.O6(CLBLM_R_X103Y112_SLICE_X163Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_AO5),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_BO5),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_AO6),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_BO6),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_CO6),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_DO6),
.Q(CLBLM_R_X103Y113_SLICE_X162Y113_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000330000)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y113_SLICE_X162Y113_CQ),
.I2(1'b1),
.I3(CLBLM_R_X103Y113_SLICE_X162Y113_A5Q),
.I4(CLBLM_R_X103Y113_SLICE_X162Y113_B5Q),
.I5(CLBLM_R_X103Y113_SLICE_X162Y113_AQ),
.O5(CLBLM_R_X103Y113_SLICE_X162Y113_DO5),
.O6(CLBLM_R_X103Y113_SLICE_X162Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303030603030)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_CLUT (
.I0(CLBLM_R_X103Y113_SLICE_X162Y113_AQ),
.I1(CLBLM_R_X103Y113_SLICE_X162Y113_CQ),
.I2(CLBLM_R_X103Y113_SLICE_X163Y113_AO6),
.I3(CLBLM_R_X103Y113_SLICE_X162Y113_A5Q),
.I4(CLBLM_R_X103Y113_SLICE_X162Y113_B5Q),
.I5(CLBLL_L_X102Y112_SLICE_X161Y112_CO6),
.O5(CLBLM_R_X103Y113_SLICE_X162Y113_CO5),
.O6(CLBLM_R_X103Y113_SLICE_X162Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffa050a050)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_BLUT (
.I0(CLBLM_R_X103Y113_SLICE_X162Y113_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X103Y113_SLICE_X163Y113_AO6),
.I3(CLBLL_L_X102Y112_SLICE_X161Y112_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X162Y113_BO5),
.O6(CLBLM_R_X103Y113_SLICE_X162Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h20d020d00020f0d0)
  ) CLBLM_R_X103Y113_SLICE_X162Y113_ALUT (
.I0(CLBLM_R_X103Y113_SLICE_X162Y113_B5Q),
.I1(CLBLL_L_X102Y112_SLICE_X161Y112_CO6),
.I2(CLBLM_R_X103Y113_SLICE_X163Y113_AO6),
.I3(CLBLM_R_X103Y113_SLICE_X162Y113_AQ),
.I4(CLBLM_R_X103Y113_SLICE_X162Y113_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X162Y113_AO5),
.O6(CLBLM_R_X103Y113_SLICE_X162Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(1'b1),
.Q(CLBLM_R_X103Y113_SLICE_X163Y113_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y113_SLICE_X163Y113_AQ),
.Q(CLBLM_R_X103Y113_SLICE_X163Y113_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y113_SLICE_X162Y113_DQ),
.Q(CLBLM_R_X103Y113_SLICE_X163Y113_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X163Y113_DO5),
.O6(CLBLM_R_X103Y113_SLICE_X163Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X163Y113_CO5),
.O6(CLBLM_R_X103Y113_SLICE_X163Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X163Y113_BO5),
.O6(CLBLM_R_X103Y113_SLICE_X163Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f0b0f030303030)
  ) CLBLM_R_X103Y113_SLICE_X163Y113_ALUT (
.I0(CLBLM_R_X103Y113_SLICE_X162Y113_DQ),
.I1(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X103Y113_SLICE_X162Y113_BQ),
.I4(CLBLM_R_X103Y113_SLICE_X163Y113_CQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y113_SLICE_X163Y113_AO5),
.O6(CLBLM_R_X103Y113_SLICE_X163Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y114_SLICE_X162Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y114_SLICE_X162Y114_AO6),
.Q(CLBLM_R_X103Y114_SLICE_X162Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y114_SLICE_X162Y114_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y114_SLICE_X162Y114_BO6),
.Q(CLBLM_R_X103Y114_SLICE_X162Y114_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y114_SLICE_X162Y114_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y114_SLICE_X162Y114_CO6),
.Q(CLBLM_R_X103Y114_SLICE_X162Y114_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X103Y114_SLICE_X162Y114_DLUT (
.I0(CLBLM_R_X103Y114_SLICE_X163Y114_AQ),
.I1(CLBLM_R_X103Y114_SLICE_X162Y114_CQ),
.I2(CLBLM_R_X103Y114_SLICE_X162Y114_AQ),
.I3(CLBLM_R_X103Y114_SLICE_X162Y114_BQ),
.I4(CLBLM_R_X103Y116_SLICE_X163Y116_B5Q),
.I5(CLBLL_L_X102Y114_SLICE_X161Y114_AQ),
.O5(CLBLM_R_X103Y114_SLICE_X162Y114_DO5),
.O6(CLBLM_R_X103Y114_SLICE_X162Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d85050cccc0000)
  ) CLBLM_R_X103Y114_SLICE_X162Y114_CLUT (
.I0(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I1(CLBLM_R_X103Y114_SLICE_X162Y114_CQ),
.I2(CLBLM_R_X103Y114_SLICE_X162Y114_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.O5(CLBLM_R_X103Y114_SLICE_X162Y114_CO5),
.O6(CLBLM_R_X103Y114_SLICE_X162Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0eac040c0eac040)
  ) CLBLM_R_X103Y114_SLICE_X162Y114_BLUT (
.I0(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I1(CLBLM_R_X103Y114_SLICE_X162Y114_BQ),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I4(CLBLM_R_X103Y114_SLICE_X163Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y114_SLICE_X162Y114_BO5),
.O6(CLBLM_R_X103Y114_SLICE_X162Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fa500000aa00)
  ) CLBLM_R_X103Y114_SLICE_X162Y114_ALUT (
.I0(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I1(1'b1),
.I2(CLBLM_R_X103Y114_SLICE_X162Y114_AQ),
.I3(CLBLM_R_X103Y115_SLICE_X162Y115_AQ),
.I4(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X103Y114_SLICE_X162Y114_AO5),
.O6(CLBLM_R_X103Y114_SLICE_X162Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y114_SLICE_X163Y114_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y114_SLICE_X163Y114_AO6),
.Q(CLBLM_R_X103Y114_SLICE_X163Y114_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y114_SLICE_X163Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y114_SLICE_X163Y114_DO5),
.O6(CLBLM_R_X103Y114_SLICE_X163Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y114_SLICE_X163Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y114_SLICE_X163Y114_CO5),
.O6(CLBLM_R_X103Y114_SLICE_X163Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7f7f7fffffffff)
  ) CLBLM_R_X103Y114_SLICE_X163Y114_BLUT (
.I0(CLBLM_R_X103Y115_SLICE_X163Y115_DQ),
.I1(CLBLM_R_X103Y115_SLICE_X163Y115_BQ),
.I2(CLBLM_R_X103Y115_SLICE_X163Y115_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X103Y115_SLICE_X163Y115_CQ),
.O5(CLBLM_R_X103Y114_SLICE_X163Y114_BO5),
.O6(CLBLM_R_X103Y114_SLICE_X163Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c03300f0f00000)
  ) CLBLM_R_X103Y114_SLICE_X163Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I2(CLBLM_R_X103Y114_SLICE_X163Y114_AQ),
.I3(CLBLM_R_X103Y116_SLICE_X163Y116_B5Q),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.O5(CLBLM_R_X103Y114_SLICE_X163Y114_AO5),
.O6(CLBLM_R_X103Y114_SLICE_X163Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y115_SLICE_X162Y115_AO5),
.Q(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y115_SLICE_X162Y115_AO6),
.Q(CLBLM_R_X103Y115_SLICE_X162Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y115_SLICE_X162Y115_BO6),
.Q(CLBLM_R_X103Y115_SLICE_X162Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y115_SLICE_X162Y115_CO6),
.Q(CLBLM_R_X103Y115_SLICE_X162Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000300000000)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y115_SLICE_X162Y115_CQ),
.I2(CLBLM_R_X103Y115_SLICE_X162Y115_AQ),
.I3(CLBLM_R_X103Y115_SLICE_X162Y115_BQ),
.I4(1'b1),
.I5(CLBLM_R_X103Y114_SLICE_X162Y114_DO6),
.O5(CLBLM_R_X103Y115_SLICE_X162Y115_DO5),
.O6(CLBLM_R_X103Y115_SLICE_X162Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ccd8cc50005000)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_CLUT (
.I0(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I1(CLBLM_R_X103Y115_SLICE_X162Y115_CQ),
.I2(CLBLM_R_X103Y115_SLICE_X162Y115_BQ),
.I3(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I4(1'b1),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X103Y115_SLICE_X162Y115_CO5),
.O6(CLBLM_R_X103Y115_SLICE_X162Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00f0f0cc00cc00)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y115_SLICE_X162Y115_BQ),
.I2(CLBLL_L_X102Y114_SLICE_X161Y114_AQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I5(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.O5(CLBLM_R_X103Y115_SLICE_X162Y115_BO5),
.O6(CLBLM_R_X103Y115_SLICE_X162Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he222f000ffffcccc)
  ) CLBLM_R_X103Y115_SLICE_X162Y115_ALUT (
.I0(CLBLM_R_X103Y114_SLICE_X162Y114_BQ),
.I1(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I2(CLBLM_R_X103Y115_SLICE_X162Y115_AQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y115_SLICE_X162Y115_AO5),
.O6(CLBLM_R_X103Y115_SLICE_X162Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y115_SLICE_X163Y115_AO6),
.Q(CLBLM_R_X103Y115_SLICE_X163Y115_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y115_SLICE_X163Y115_BO6),
.Q(CLBLM_R_X103Y115_SLICE_X163Y115_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y115_SLICE_X163Y115_CO6),
.Q(CLBLM_R_X103Y115_SLICE_X163Y115_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y115_SLICE_X163Y115_DO6),
.Q(CLBLM_R_X103Y115_SLICE_X163Y115_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8cc00cc00cc00cc0)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_DLUT (
.I0(CLBLM_R_X103Y115_SLICE_X163Y115_BQ),
.I1(CLBLM_R_X103Y113_SLICE_X163Y113_AO5),
.I2(CLBLM_R_X103Y115_SLICE_X163Y115_DQ),
.I3(CLBLM_R_X103Y116_SLICE_X163Y116_CO6),
.I4(CLBLM_R_X103Y115_SLICE_X163Y115_CQ),
.I5(CLBLM_R_X103Y115_SLICE_X163Y115_AQ),
.O5(CLBLM_R_X103Y115_SLICE_X163Y115_DO5),
.O6(CLBLM_R_X103Y115_SLICE_X163Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8cccc0000cccc000)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_CLUT (
.I0(CLBLM_R_X103Y115_SLICE_X163Y115_BQ),
.I1(CLBLM_R_X103Y113_SLICE_X163Y113_AO5),
.I2(CLBLM_R_X103Y115_SLICE_X163Y115_DQ),
.I3(CLBLM_R_X103Y116_SLICE_X163Y116_CO6),
.I4(CLBLM_R_X103Y115_SLICE_X163Y115_CQ),
.I5(CLBLM_R_X103Y115_SLICE_X163Y115_AQ),
.O5(CLBLM_R_X103Y115_SLICE_X163Y115_CO5),
.O6(CLBLM_R_X103Y115_SLICE_X163Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he6cc0000cccc0000)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_BLUT (
.I0(CLBLM_R_X103Y115_SLICE_X163Y115_CQ),
.I1(CLBLM_R_X103Y115_SLICE_X163Y115_BQ),
.I2(CLBLM_R_X103Y115_SLICE_X163Y115_AQ),
.I3(CLBLM_R_X103Y115_SLICE_X163Y115_DQ),
.I4(CLBLM_R_X103Y113_SLICE_X163Y113_AO5),
.I5(CLBLM_R_X103Y116_SLICE_X163Y116_CO6),
.O5(CLBLM_R_X103Y115_SLICE_X163Y115_BO5),
.O6(CLBLM_R_X103Y115_SLICE_X163Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f00000f0f00000)
  ) CLBLM_R_X103Y115_SLICE_X163Y115_ALUT (
.I0(CLBLM_R_X103Y115_SLICE_X163Y115_CQ),
.I1(CLBLM_R_X103Y115_SLICE_X163Y115_BQ),
.I2(CLBLM_R_X103Y115_SLICE_X163Y115_AQ),
.I3(CLBLM_R_X103Y115_SLICE_X163Y115_DQ),
.I4(CLBLM_R_X103Y113_SLICE_X163Y113_AO5),
.I5(CLBLM_R_X103Y116_SLICE_X163Y116_CO6),
.O5(CLBLM_R_X103Y115_SLICE_X163Y115_AO5),
.O6(CLBLM_R_X103Y115_SLICE_X163Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y117_SLICE_X162Y117_BO6),
.Q(CLBLM_R_X103Y116_SLICE_X162Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y116_SLICE_X163Y116_DQ),
.Q(CLBLM_R_X103Y116_SLICE_X162Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y116_SLICE_X162Y116_AO6),
.Q(CLBLM_R_X103Y116_SLICE_X162Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y116_SLICE_X162Y116_BO6),
.Q(CLBLM_R_X103Y116_SLICE_X162Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y116_SLICE_X162Y116_CO6),
.Q(CLBLM_R_X103Y116_SLICE_X162Y116_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a00aa00ffffffff)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_DLUT (
.I0(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I1(1'b1),
.I2(CLBLM_R_X103Y116_SLICE_X163Y116_DQ),
.I3(CLBLM_R_X103Y116_SLICE_X162Y116_A5Q),
.I4(CLBLM_R_X103Y116_SLICE_X162Y116_B5Q),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X103Y116_SLICE_X162Y116_DO5),
.O6(CLBLM_R_X103Y116_SLICE_X162Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc00003333)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y116_SLICE_X162Y116_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X103Y116_SLICE_X162Y116_DO6),
.I5(CLBLM_R_X103Y117_SLICE_X162Y117_BO6),
.O5(CLBLM_R_X103Y116_SLICE_X162Y116_CO5),
.O6(CLBLM_R_X103Y116_SLICE_X162Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00f0f0cc00cc00)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y116_SLICE_X162Y116_BQ),
.I2(CLBLM_R_X103Y116_SLICE_X162Y116_AQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I5(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.O5(CLBLM_R_X103Y116_SLICE_X162Y116_BO5),
.O6(CLBLM_R_X103Y116_SLICE_X162Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000b888f000b888)
  ) CLBLM_R_X103Y116_SLICE_X162Y116_ALUT (
.I0(CLBLL_L_X102Y115_SLICE_X161Y115_AQ),
.I1(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I2(CLBLM_R_X103Y116_SLICE_X162Y116_AQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y116_SLICE_X162Y116_AO5),
.O6(CLBLM_R_X103Y116_SLICE_X162Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y116_SLICE_X163Y116_AO5),
.Q(CLBLM_R_X103Y116_SLICE_X163Y116_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y116_SLICE_X163Y116_CO5),
.Q(CLBLM_R_X103Y116_SLICE_X163Y116_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y116_SLICE_X163Y116_AO6),
.Q(CLBLM_R_X103Y116_SLICE_X163Y116_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y116_SLICE_X163Y116_BO6),
.Q(CLBLM_R_X103Y116_SLICE_X163Y116_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y116_SLICE_X163Y116_DO6),
.Q(CLBLM_R_X103Y116_SLICE_X163Y116_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000003)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X103Y116_SLICE_X163Y116_BQ),
.I2(CLBLM_R_X103Y116_SLICE_X163Y116_A5Q),
.I3(CLBLM_R_X103Y116_SLICE_X162Y116_CQ),
.I4(CLBLM_R_X103Y116_SLICE_X163Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y116_SLICE_X163Y116_DO5),
.O6(CLBLM_R_X103Y116_SLICE_X163Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444444fb404040)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_CLUT (
.I0(CLBLM_R_X103Y113_SLICE_X163Y113_BQ),
.I1(CLBLM_R_X103Y115_SLICE_X162Y115_A5Q),
.I2(CLBLM_R_X103Y117_SLICE_X162Y117_CO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X103Y116_SLICE_X163Y116_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y116_SLICE_X163Y116_CO5),
.O6(CLBLM_R_X103Y116_SLICE_X163Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111111111111211)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_BLUT (
.I0(CLBLM_R_X103Y116_SLICE_X163Y116_BQ),
.I1(CLBLM_R_X103Y116_SLICE_X162Y116_DO6),
.I2(CLBLM_R_X103Y116_SLICE_X163Y116_AQ),
.I3(CLBLM_R_X103Y117_SLICE_X162Y117_BO6),
.I4(CLBLM_R_X103Y116_SLICE_X162Y116_CQ),
.I5(CLBLM_R_X103Y116_SLICE_X163Y116_A5Q),
.O5(CLBLM_R_X103Y116_SLICE_X163Y116_BO5),
.O6(CLBLM_R_X103Y116_SLICE_X163Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111221103031203)
  ) CLBLM_R_X103Y116_SLICE_X163Y116_ALUT (
.I0(CLBLM_R_X103Y116_SLICE_X163Y116_AQ),
.I1(CLBLM_R_X103Y116_SLICE_X162Y116_DO6),
.I2(CLBLM_R_X103Y116_SLICE_X163Y116_A5Q),
.I3(CLBLM_R_X103Y117_SLICE_X162Y117_BO6),
.I4(CLBLM_R_X103Y116_SLICE_X162Y116_CQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y116_SLICE_X163Y116_AO5),
.O6(CLBLM_R_X103Y116_SLICE_X163Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y117_SLICE_X162Y117_AO6),
.Q(CLBLM_R_X103Y117_SLICE_X162Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y117_SLICE_X162Y117_DO5),
.O6(CLBLM_R_X103Y117_SLICE_X162Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500ae00ae)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_CLUT (
.I0(CLBLM_R_X103Y116_SLICE_X162Y116_AQ),
.I1(CLBLM_R_X103Y115_SLICE_X162Y115_DO6),
.I2(CLBLL_L_X102Y115_SLICE_X161Y115_DO6),
.I3(CLBLM_R_X103Y114_SLICE_X163Y114_BO6),
.I4(1'b1),
.I5(CLBLM_R_X103Y116_SLICE_X162Y116_BQ),
.O5(CLBLM_R_X103Y117_SLICE_X162Y117_CO5),
.O6(CLBLM_R_X103Y117_SLICE_X162Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00004cc400004ccc)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_BLUT (
.I0(CLBLM_R_X103Y115_SLICE_X162Y115_DO6),
.I1(CLBLM_R_X103Y116_SLICE_X163Y116_CO6),
.I2(CLBLM_R_X103Y116_SLICE_X162Y116_AQ),
.I3(CLBLM_R_X103Y116_SLICE_X162Y116_BQ),
.I4(CLBLM_R_X103Y114_SLICE_X163Y114_BO6),
.I5(CLBLL_L_X102Y115_SLICE_X161Y115_DO6),
.O5(CLBLM_R_X103Y117_SLICE_X162Y117_BO5),
.O6(CLBLM_R_X103Y117_SLICE_X162Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0e00000f0c0000)
  ) CLBLM_R_X103Y117_SLICE_X162Y117_ALUT (
.I0(CLBLM_R_X103Y118_SLICE_X162Y118_B5Q),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(CLBLM_R_X103Y117_SLICE_X162Y117_AQ),
.I3(CLBLM_R_X103Y118_SLICE_X163Y118_BQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X103Y117_SLICE_X163Y117_DQ),
.O5(CLBLM_R_X103Y117_SLICE_X162Y117_AO5),
.O6(CLBLM_R_X103Y117_SLICE_X162Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y117_SLICE_X163Y117_AO6),
.Q(CLBLM_R_X103Y117_SLICE_X163Y117_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y117_SLICE_X163Y117_BO6),
.Q(CLBLM_R_X103Y117_SLICE_X163Y117_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_C_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y117_SLICE_X163Y117_CO6),
.Q(CLBLM_R_X103Y117_SLICE_X163Y117_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_D_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y117_SLICE_X163Y117_DO6),
.Q(CLBLM_R_X103Y117_SLICE_X163Y117_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000100010001)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_DLUT (
.I0(CLBLM_R_X103Y117_SLICE_X162Y117_AQ),
.I1(CLBLM_R_X103Y117_SLICE_X163Y117_CQ),
.I2(CLBLM_R_X103Y117_SLICE_X163Y117_BQ),
.I3(CLBLM_R_X103Y117_SLICE_X163Y117_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y117_SLICE_X163Y117_DO5),
.O6(CLBLM_R_X103Y117_SLICE_X163Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222222202200)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_R_X103Y117_SLICE_X163Y117_CQ),
.I2(CLBLM_R_X103Y117_SLICE_X163Y117_DQ),
.I3(CLBLM_R_X103Y118_SLICE_X163Y118_BQ),
.I4(CLBLM_R_X103Y118_SLICE_X162Y118_B5Q),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLM_R_X103Y117_SLICE_X163Y117_CO5),
.O6(CLBLM_R_X103Y117_SLICE_X163Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030302030303000)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_BLUT (
.I0(CLBLM_R_X103Y118_SLICE_X162Y118_B5Q),
.I1(CLBLM_R_X103Y117_SLICE_X163Y117_BQ),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X103Y118_SLICE_X163Y118_BQ),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLM_R_X103Y117_SLICE_X163Y117_DQ),
.O5(CLBLM_R_X103Y117_SLICE_X163Y117_BO5),
.O6(CLBLM_R_X103Y117_SLICE_X163Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f080)
  ) CLBLM_R_X103Y117_SLICE_X163Y117_ALUT (
.I0(CLBLM_R_X103Y118_SLICE_X162Y118_B5Q),
.I1(CLBLM_R_X103Y117_SLICE_X163Y117_DQ),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X103Y118_SLICE_X163Y118_BQ),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLM_R_X103Y117_SLICE_X163Y117_AQ),
.O5(CLBLM_R_X103Y117_SLICE_X163Y117_AO5),
.O6(CLBLM_R_X103Y117_SLICE_X163Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y118_SLICE_X162Y118_A5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y118_SLICE_X162Y118_AO5),
.Q(CLBLM_R_X103Y118_SLICE_X162Y118_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y118_SLICE_X162Y118_B5_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y117_SLICE_X163Y117_DQ),
.Q(CLBLM_R_X103Y118_SLICE_X162Y118_B5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y118_SLICE_X162Y118_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y118_SLICE_X162Y118_AO6),
.Q(CLBLM_R_X103Y118_SLICE_X162Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y118_SLICE_X162Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y118_SLICE_X162Y118_BO6),
.Q(CLBLM_R_X103Y118_SLICE_X162Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y118_SLICE_X162Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y118_SLICE_X162Y118_DO5),
.O6(CLBLM_R_X103Y118_SLICE_X162Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a8a88888)
  ) CLBLM_R_X103Y118_SLICE_X162Y118_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y113_IOB_X1Y114_I),
.I2(CLBLM_R_X103Y117_SLICE_X163Y117_DQ),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I4(CLBLM_R_X103Y118_SLICE_X162Y118_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X103Y118_SLICE_X162Y118_CO5),
.O6(CLBLM_R_X103Y118_SLICE_X162Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a000000aa000000)
  ) CLBLM_R_X103Y118_SLICE_X162Y118_BLUT (
.I0(CLBLM_R_X103Y118_SLICE_X162Y118_BQ),
.I1(CLBLM_R_X103Y112_SLICE_X162Y112_A5Q),
.I2(CLBLM_R_X103Y118_SLICE_X162Y118_AQ),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X103Y118_SLICE_X162Y118_A5Q),
.O5(CLBLM_R_X103Y118_SLICE_X162Y118_BO5),
.O6(CLBLM_R_X103Y118_SLICE_X162Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c0000006a000000)
  ) CLBLM_R_X103Y118_SLICE_X162Y118_ALUT (
.I0(CLBLM_R_X103Y118_SLICE_X162Y118_A5Q),
.I1(CLBLM_R_X103Y112_SLICE_X162Y112_A5Q),
.I2(CLBLM_R_X103Y118_SLICE_X162Y118_AQ),
.I3(CLBLL_L_X102Y115_SLICE_X161Y115_A5Q),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y118_SLICE_X162Y118_AO5),
.O6(CLBLM_R_X103Y118_SLICE_X162Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDPE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y118_SLICE_X163Y118_A_FDPE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_R_X103Y118_SLICE_X162Y118_CO5),
.PRE(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.Q(CLBLM_R_X103Y118_SLICE_X163Y118_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y118_SLICE_X163Y118_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y118_SLICE_X163Y118_AQ),
.Q(CLBLM_R_X103Y118_SLICE_X163Y118_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y118_SLICE_X163Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y118_SLICE_X163Y118_DO5),
.O6(CLBLM_R_X103Y118_SLICE_X163Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y118_SLICE_X163Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y118_SLICE_X163Y118_CO5),
.O6(CLBLM_R_X103Y118_SLICE_X163Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y118_SLICE_X163Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y118_SLICE_X163Y118_BO5),
.O6(CLBLM_R_X103Y118_SLICE_X163Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y118_SLICE_X163Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y118_SLICE_X163Y118_AO5),
.O6(CLBLM_R_X103Y118_SLICE_X163Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y119_SLICE_X162Y119_AO6),
.Q(CLBLM_R_X103Y119_SLICE_X162Y119_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_B_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y119_SLICE_X162Y119_BO6),
.Q(CLBLM_R_X103Y119_SLICE_X162Y119_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555ffffffff)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_DLUT (
.I0(CLBLM_R_X103Y118_SLICE_X162Y118_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X103Y112_SLICE_X162Y112_A5Q),
.O5(CLBLM_R_X103Y119_SLICE_X162Y119_DO5),
.O6(CLBLM_R_X103Y119_SLICE_X162Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_CLUT (
.I0(CLBLM_R_X103Y118_SLICE_X162Y118_A5Q),
.I1(CLBLM_R_X103Y118_SLICE_X162Y118_AQ),
.I2(CLBLM_R_X103Y119_SLICE_X162Y119_AQ),
.I3(CLBLM_R_X103Y112_SLICE_X162Y112_A5Q),
.I4(CLBLM_R_X103Y119_SLICE_X162Y119_BQ),
.I5(CLBLM_R_X103Y118_SLICE_X162Y118_BQ),
.O5(CLBLM_R_X103Y119_SLICE_X162Y119_CO5),
.O6(CLBLM_R_X103Y119_SLICE_X162Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8828888888888888)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_BLUT (
.I0(CLBLM_R_X103Y118_SLICE_X162Y118_CO6),
.I1(CLBLM_R_X103Y119_SLICE_X162Y119_BQ),
.I2(CLBLM_R_X103Y118_SLICE_X162Y118_A5Q),
.I3(CLBLM_R_X103Y119_SLICE_X162Y119_DO6),
.I4(CLBLM_R_X103Y118_SLICE_X162Y118_BQ),
.I5(CLBLM_R_X103Y119_SLICE_X162Y119_AQ),
.O5(CLBLM_R_X103Y119_SLICE_X162Y119_BO5),
.O6(CLBLM_R_X103Y119_SLICE_X162Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2aaaaaaa80000000)
  ) CLBLM_R_X103Y119_SLICE_X162Y119_ALUT (
.I0(CLBLM_R_X103Y118_SLICE_X162Y118_CO6),
.I1(CLBLM_R_X103Y118_SLICE_X162Y118_BQ),
.I2(CLBLM_R_X103Y118_SLICE_X162Y118_AQ),
.I3(CLBLM_R_X103Y112_SLICE_X162Y112_A5Q),
.I4(CLBLM_R_X103Y118_SLICE_X162Y118_A5Q),
.I5(CLBLM_R_X103Y119_SLICE_X162Y119_AQ),
.O5(CLBLM_R_X103Y119_SLICE_X162Y119_AO5),
.O6(CLBLM_R_X103Y119_SLICE_X162Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y119_SLICE_X163Y119_DO5),
.O6(CLBLM_R_X103Y119_SLICE_X163Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y119_SLICE_X163Y119_CO5),
.O6(CLBLM_R_X103Y119_SLICE_X163Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y119_SLICE_X163Y119_BO5),
.O6(CLBLM_R_X103Y119_SLICE_X163Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y119_SLICE_X163Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y119_SLICE_X163Y119_AO5),
.O6(CLBLM_R_X103Y119_SLICE_X163Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_DO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_CO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_BO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X162Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X162Y122_AO5),
.O6(CLBLM_R_X103Y122_SLICE_X162Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_A_FDCE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.CLR(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.D(CLBLM_R_X103Y122_SLICE_X163Y122_AO6),
.Q(CLBLM_R_X103Y122_SLICE_X163Y122_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_DO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_CO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_BO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X103Y122_SLICE_X163Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X103Y122_SLICE_X163Y122_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y122_SLICE_X163Y122_AO5),
.O6(CLBLM_R_X103Y122_SLICE_X163Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X102Y107_SLICE_X160Y107_AQ),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X102Y107_SLICE_X160Y107_A5Q),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X102Y107_SLICE_X160Y107_BQ),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_I),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLM_R_X103Y108_SLICE_X162Y108_CO6),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLM_R_X103Y109_SLICE_X163Y109_AO5),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(1'b1),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(1'b0),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(1'b0),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(1'b0),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(1'b0),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(1'b1),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(1'b0),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(1'b0),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(1'b0),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(1'b0),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(1'b0),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(1'b0),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(1'b0),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(1'b0),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(1'b0),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(1'b0),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(1'b0),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(1'b0),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(1'b0),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(1'b0),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(1'b0),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(1'b0),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(1'b0),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(1'b0),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(1'b0),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(1'b0),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(1'b0),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(1'b0),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(1'b0),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(1'b0),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(1'b0),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(1'b1),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(1'b0),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLM_R_X103Y119_SLICE_X162Y119_BQ),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(1'b0),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(1'b1),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y115_OBUF (
.I(1'b1),
.O(RIOB33_X105Y115_IOB_X1Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y115_IOB_X1Y116_OBUF (
.I(1'b1),
.O(RIOB33_X105Y115_IOB_X1Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y117_OBUF (
.I(1'b1),
.O(RIOB33_X105Y117_IOB_X1Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y117_IOB_X1Y118_OBUF (
.I(1'b1),
.O(RIOB33_X105Y117_IOB_X1Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y119_OBUF (
.I(1'b1),
.O(RIOB33_X105Y119_IOB_X1Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y119_IOB_X1Y120_OBUF (
.I(1'b1),
.O(RIOB33_X105Y119_IOB_X1Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y121_OBUF (
.I(1'b1),
.O(RIOB33_X105Y121_IOB_X1Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y121_IOB_X1Y122_OBUF (
.I(1'b1),
.O(RIOB33_X105Y121_IOB_X1Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y123_OBUF (
.I(CLBLM_R_X103Y122_SLICE_X163Y122_AQ),
.O(RIOB33_X105Y123_IOB_X1Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y123_IOB_X1Y124_OBUF (
.I(1'b1),
.O(RIOB33_X105Y123_IOB_X1Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y125_OBUF (
.I(1'b0),
.O(RIOB33_X105Y125_IOB_X1Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y125_IOB_X1Y126_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y125_IOB_X1Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y127_IOB_X1Y127_OBUF (
.I(1'b0),
.O(RIOB33_X105Y127_IOB_X1Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y129_OBUF (
.I(1'b0),
.O(RIOB33_X105Y129_IOB_X1Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y129_IOB_X1Y130_OBUF (
.I(1'b0),
.O(RIOB33_X105Y129_IOB_X1Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y131_OBUF (
.I(1'b0),
.O(RIOB33_X105Y131_IOB_X1Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y131_IOB_X1Y132_OBUF (
.I(1'b0),
.O(RIOB33_X105Y131_IOB_X1Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y133_OBUF (
.I(1'b0),
.O(RIOB33_X105Y133_IOB_X1Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y133_IOB_X1Y134_OBUF (
.I(1'b0),
.O(RIOB33_X105Y133_IOB_X1Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y135_OBUF (
.I(1'b0),
.O(RIOB33_X105Y135_IOB_X1Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y135_IOB_X1Y136_OBUF (
.I(1'b0),
.O(RIOB33_X105Y135_IOB_X1Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y137_OBUF (
.I(1'b0),
.O(RIOB33_X105Y137_IOB_X1Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y137_IOB_X1Y138_OBUF (
.I(1'b0),
.O(RIOB33_X105Y137_IOB_X1Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y139_OBUF (
.I(1'b0),
.O(RIOB33_X105Y139_IOB_X1Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y139_IOB_X1Y140_OBUF (
.I(CLBLL_L_X102Y107_SLICE_X160Y107_CQ),
.O(RIOB33_X105Y139_IOB_X1Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y141_OBUF (
.I(CLBLM_R_X103Y117_SLICE_X163Y117_DQ),
.O(RIOB33_X105Y141_IOB_X1Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y141_IOB_X1Y142_OBUF (
.I(CLBLM_R_X103Y113_SLICE_X162Y113_DQ),
.O(RIOB33_X105Y141_IOB_X1Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y143_OBUF (
.I(CLBLM_R_X103Y116_SLICE_X163Y116_DQ),
.O(RIOB33_X105Y143_IOB_X1Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y143_IOB_X1Y144_OBUF (
.I(1'b0),
.O(RIOB33_X105Y143_IOB_X1Y144_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y145_OBUF (
.I(CLBLM_R_X103Y112_SLICE_X162Y112_A5Q),
.O(RIOB33_X105Y145_IOB_X1Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y145_IOB_X1Y146_OBUF (
.I(CLBLM_R_X103Y118_SLICE_X162Y118_AQ),
.O(RIOB33_X105Y145_IOB_X1Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y147_OBUF (
.I(CLBLM_R_X103Y118_SLICE_X162Y118_A5Q),
.O(RIOB33_X105Y147_IOB_X1Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y147_IOB_X1Y148_OBUF (
.I(CLBLM_R_X103Y118_SLICE_X162Y118_BQ),
.O(RIOB33_X105Y147_IOB_X1Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y149_IOB_X1Y149_OBUF (
.I(CLBLM_R_X103Y119_SLICE_X162Y119_AQ),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_OPAD)
  );
  assign CLBLL_L_X102Y107_SLICE_X160Y107_A = CLBLL_L_X102Y107_SLICE_X160Y107_AO6;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_B = CLBLL_L_X102Y107_SLICE_X160Y107_BO6;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_C = CLBLL_L_X102Y107_SLICE_X160Y107_CO6;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_D = CLBLL_L_X102Y107_SLICE_X160Y107_DO6;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_AMUX = CLBLL_L_X102Y107_SLICE_X160Y107_A5Q;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_A = CLBLL_L_X102Y107_SLICE_X161Y107_AO6;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_B = CLBLL_L_X102Y107_SLICE_X161Y107_BO6;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_C = CLBLL_L_X102Y107_SLICE_X161Y107_CO6;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_D = CLBLL_L_X102Y107_SLICE_X161Y107_DO6;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_A = CLBLL_L_X102Y108_SLICE_X160Y108_AO6;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_B = CLBLL_L_X102Y108_SLICE_X160Y108_BO6;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_C = CLBLL_L_X102Y108_SLICE_X160Y108_CO6;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_D = CLBLL_L_X102Y108_SLICE_X160Y108_DO6;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_A = CLBLL_L_X102Y108_SLICE_X161Y108_AO6;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_B = CLBLL_L_X102Y108_SLICE_X161Y108_BO6;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_C = CLBLL_L_X102Y108_SLICE_X161Y108_CO6;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_D = CLBLL_L_X102Y108_SLICE_X161Y108_DO6;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_BMUX = CLBLL_L_X102Y108_SLICE_X161Y108_B5Q;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_A = CLBLL_L_X102Y109_SLICE_X160Y109_AO6;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_B = CLBLL_L_X102Y109_SLICE_X160Y109_BO6;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_C = CLBLL_L_X102Y109_SLICE_X160Y109_CO6;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_D = CLBLL_L_X102Y109_SLICE_X160Y109_DO6;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_AMUX = CLBLL_L_X102Y109_SLICE_X160Y109_A5Q;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_BMUX = CLBLL_L_X102Y109_SLICE_X160Y109_B5Q;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_CMUX = CLBLL_L_X102Y109_SLICE_X160Y109_C5Q;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_A = CLBLL_L_X102Y109_SLICE_X161Y109_AO6;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_B = CLBLL_L_X102Y109_SLICE_X161Y109_BO6;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_C = CLBLL_L_X102Y109_SLICE_X161Y109_CO6;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_D = CLBLL_L_X102Y109_SLICE_X161Y109_DO6;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_AMUX = CLBLL_L_X102Y109_SLICE_X161Y109_AO5;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_BMUX = CLBLL_L_X102Y109_SLICE_X161Y109_B5Q;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_CMUX = CLBLL_L_X102Y109_SLICE_X161Y109_CO5;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_A = CLBLL_L_X102Y110_SLICE_X160Y110_AO6;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_B = CLBLL_L_X102Y110_SLICE_X160Y110_BO6;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_C = CLBLL_L_X102Y110_SLICE_X160Y110_CO6;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_D = CLBLL_L_X102Y110_SLICE_X160Y110_DO6;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_AMUX = CLBLL_L_X102Y110_SLICE_X160Y110_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_BMUX = CLBLL_L_X102Y110_SLICE_X160Y110_B5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_CMUX = CLBLL_L_X102Y110_SLICE_X160Y110_C5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_DMUX = CLBLL_L_X102Y110_SLICE_X160Y110_D5Q;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_A = CLBLL_L_X102Y110_SLICE_X161Y110_AO6;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_B = CLBLL_L_X102Y110_SLICE_X161Y110_BO6;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_C = CLBLL_L_X102Y110_SLICE_X161Y110_CO6;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_D = CLBLL_L_X102Y110_SLICE_X161Y110_DO6;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_AMUX = CLBLL_L_X102Y110_SLICE_X161Y110_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_BMUX = CLBLL_L_X102Y110_SLICE_X161Y110_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A = CLBLL_L_X102Y111_SLICE_X160Y111_AO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B = CLBLL_L_X102Y111_SLICE_X160Y111_BO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C = CLBLL_L_X102Y111_SLICE_X160Y111_CO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D = CLBLL_L_X102Y111_SLICE_X160Y111_DO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_AMUX = CLBLL_L_X102Y111_SLICE_X160Y111_A5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_BMUX = CLBLL_L_X102Y111_SLICE_X160Y111_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_CMUX = CLBLL_L_X102Y111_SLICE_X160Y111_C5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A = CLBLL_L_X102Y111_SLICE_X161Y111_AO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B = CLBLL_L_X102Y111_SLICE_X161Y111_BO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C = CLBLL_L_X102Y111_SLICE_X161Y111_CO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D = CLBLL_L_X102Y111_SLICE_X161Y111_DO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A = CLBLL_L_X102Y112_SLICE_X160Y112_AO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B = CLBLL_L_X102Y112_SLICE_X160Y112_BO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C = CLBLL_L_X102Y112_SLICE_X160Y112_CO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D = CLBLL_L_X102Y112_SLICE_X160Y112_DO6;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_AMUX = CLBLL_L_X102Y112_SLICE_X160Y112_A5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_BMUX = CLBLL_L_X102Y112_SLICE_X160Y112_B5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_CMUX = CLBLL_L_X102Y112_SLICE_X160Y112_C5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A = CLBLL_L_X102Y112_SLICE_X161Y112_AO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B = CLBLL_L_X102Y112_SLICE_X161Y112_BO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C = CLBLL_L_X102Y112_SLICE_X161Y112_CO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D = CLBLL_L_X102Y112_SLICE_X161Y112_DO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_AMUX = CLBLL_L_X102Y112_SLICE_X161Y112_A5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_BMUX = CLBLL_L_X102Y112_SLICE_X161Y112_B5Q;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A = CLBLL_L_X102Y113_SLICE_X160Y113_AO6;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B = CLBLL_L_X102Y113_SLICE_X160Y113_BO6;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C = CLBLL_L_X102Y113_SLICE_X160Y113_CO6;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D = CLBLL_L_X102Y113_SLICE_X160Y113_DO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A = CLBLL_L_X102Y113_SLICE_X161Y113_AO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B = CLBLL_L_X102Y113_SLICE_X161Y113_BO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C = CLBLL_L_X102Y113_SLICE_X161Y113_CO6;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D = CLBLL_L_X102Y113_SLICE_X161Y113_DO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A = CLBLL_L_X102Y114_SLICE_X160Y114_AO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B = CLBLL_L_X102Y114_SLICE_X160Y114_BO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C = CLBLL_L_X102Y114_SLICE_X160Y114_CO6;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D = CLBLL_L_X102Y114_SLICE_X160Y114_DO6;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A = CLBLL_L_X102Y114_SLICE_X161Y114_AO6;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B = CLBLL_L_X102Y114_SLICE_X161Y114_BO6;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C = CLBLL_L_X102Y114_SLICE_X161Y114_CO6;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D = CLBLL_L_X102Y114_SLICE_X161Y114_DO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A = CLBLL_L_X102Y115_SLICE_X160Y115_AO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B = CLBLL_L_X102Y115_SLICE_X160Y115_BO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C = CLBLL_L_X102Y115_SLICE_X160Y115_CO6;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D = CLBLL_L_X102Y115_SLICE_X160Y115_DO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A = CLBLL_L_X102Y115_SLICE_X161Y115_AO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B = CLBLL_L_X102Y115_SLICE_X161Y115_BO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C = CLBLL_L_X102Y115_SLICE_X161Y115_CO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D = CLBLL_L_X102Y115_SLICE_X161Y115_DO6;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_AMUX = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A = CLBLM_R_X103Y108_SLICE_X162Y108_AO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B = CLBLM_R_X103Y108_SLICE_X162Y108_BO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C = CLBLM_R_X103Y108_SLICE_X162Y108_CO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D = CLBLM_R_X103Y108_SLICE_X162Y108_DO6;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_AMUX = CLBLM_R_X103Y108_SLICE_X162Y108_A5Q;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_BMUX = CLBLM_R_X103Y108_SLICE_X162Y108_B5Q;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_CMUX = CLBLM_R_X103Y108_SLICE_X162Y108_CO5;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A = CLBLM_R_X103Y108_SLICE_X163Y108_AO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B = CLBLM_R_X103Y108_SLICE_X163Y108_BO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C = CLBLM_R_X103Y108_SLICE_X163Y108_CO6;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D = CLBLM_R_X103Y108_SLICE_X163Y108_DO6;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_A = CLBLM_R_X103Y109_SLICE_X162Y109_AO6;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_B = CLBLM_R_X103Y109_SLICE_X162Y109_BO6;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_C = CLBLM_R_X103Y109_SLICE_X162Y109_CO6;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_D = CLBLM_R_X103Y109_SLICE_X162Y109_DO6;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_AMUX = CLBLM_R_X103Y109_SLICE_X162Y109_A5Q;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_BMUX = CLBLM_R_X103Y109_SLICE_X162Y109_B5Q;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_CMUX = CLBLM_R_X103Y109_SLICE_X162Y109_CO5;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_A = CLBLM_R_X103Y109_SLICE_X163Y109_AO6;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_B = CLBLM_R_X103Y109_SLICE_X163Y109_BO6;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_C = CLBLM_R_X103Y109_SLICE_X163Y109_CO6;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_D = CLBLM_R_X103Y109_SLICE_X163Y109_DO6;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_AMUX = CLBLM_R_X103Y109_SLICE_X163Y109_AO5;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_BMUX = CLBLM_R_X103Y109_SLICE_X163Y109_B5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_A = CLBLM_R_X103Y110_SLICE_X162Y110_AO6;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_B = CLBLM_R_X103Y110_SLICE_X162Y110_BO6;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_C = CLBLM_R_X103Y110_SLICE_X162Y110_CO6;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_D = CLBLM_R_X103Y110_SLICE_X162Y110_DO6;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_AMUX = CLBLM_R_X103Y110_SLICE_X162Y110_A5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_BMUX = CLBLM_R_X103Y110_SLICE_X162Y110_B5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_CMUX = CLBLM_R_X103Y110_SLICE_X162Y110_C5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_DMUX = CLBLM_R_X103Y110_SLICE_X162Y110_D5Q;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_A = CLBLM_R_X103Y110_SLICE_X163Y110_AO6;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_B = CLBLM_R_X103Y110_SLICE_X163Y110_BO6;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_C = CLBLM_R_X103Y110_SLICE_X163Y110_CO6;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_D = CLBLM_R_X103Y110_SLICE_X163Y110_DO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A = CLBLM_R_X103Y111_SLICE_X162Y111_AO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B = CLBLM_R_X103Y111_SLICE_X162Y111_BO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C = CLBLM_R_X103Y111_SLICE_X162Y111_CO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D = CLBLM_R_X103Y111_SLICE_X162Y111_DO6;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_AMUX = CLBLM_R_X103Y111_SLICE_X162Y111_A5Q;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_BMUX = CLBLM_R_X103Y111_SLICE_X162Y111_B5Q;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A = CLBLM_R_X103Y111_SLICE_X163Y111_AO6;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B = CLBLM_R_X103Y111_SLICE_X163Y111_BO6;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C = CLBLM_R_X103Y111_SLICE_X163Y111_CO6;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D = CLBLM_R_X103Y111_SLICE_X163Y111_DO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A = CLBLM_R_X103Y112_SLICE_X162Y112_AO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B = CLBLM_R_X103Y112_SLICE_X162Y112_BO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C = CLBLM_R_X103Y112_SLICE_X162Y112_CO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D = CLBLM_R_X103Y112_SLICE_X162Y112_DO6;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_AMUX = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A = CLBLM_R_X103Y112_SLICE_X163Y112_AO6;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B = CLBLM_R_X103Y112_SLICE_X163Y112_BO6;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C = CLBLM_R_X103Y112_SLICE_X163Y112_CO6;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D = CLBLM_R_X103Y112_SLICE_X163Y112_DO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A = CLBLM_R_X103Y113_SLICE_X162Y113_AO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B = CLBLM_R_X103Y113_SLICE_X162Y113_BO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C = CLBLM_R_X103Y113_SLICE_X162Y113_CO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D = CLBLM_R_X103Y113_SLICE_X162Y113_DO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_AMUX = CLBLM_R_X103Y113_SLICE_X162Y113_A5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_BMUX = CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A = CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B = CLBLM_R_X103Y113_SLICE_X163Y113_BO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C = CLBLM_R_X103Y113_SLICE_X163Y113_CO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D = CLBLM_R_X103Y113_SLICE_X163Y113_DO6;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_AMUX = CLBLM_R_X103Y113_SLICE_X163Y113_AO5;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_A = CLBLM_R_X103Y114_SLICE_X162Y114_AO6;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_B = CLBLM_R_X103Y114_SLICE_X162Y114_BO6;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_C = CLBLM_R_X103Y114_SLICE_X162Y114_CO6;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_D = CLBLM_R_X103Y114_SLICE_X162Y114_DO6;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_A = CLBLM_R_X103Y114_SLICE_X163Y114_AO6;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_B = CLBLM_R_X103Y114_SLICE_X163Y114_BO6;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_C = CLBLM_R_X103Y114_SLICE_X163Y114_CO6;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_D = CLBLM_R_X103Y114_SLICE_X163Y114_DO6;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A = CLBLM_R_X103Y115_SLICE_X162Y115_AO6;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B = CLBLM_R_X103Y115_SLICE_X162Y115_BO6;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C = CLBLM_R_X103Y115_SLICE_X162Y115_CO6;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D = CLBLM_R_X103Y115_SLICE_X162Y115_DO6;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_AMUX = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A = CLBLM_R_X103Y115_SLICE_X163Y115_AO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B = CLBLM_R_X103Y115_SLICE_X163Y115_BO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C = CLBLM_R_X103Y115_SLICE_X163Y115_CO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D = CLBLM_R_X103Y115_SLICE_X163Y115_DO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A = CLBLM_R_X103Y116_SLICE_X162Y116_AO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B = CLBLM_R_X103Y116_SLICE_X162Y116_BO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C = CLBLM_R_X103Y116_SLICE_X162Y116_CO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D = CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_AMUX = CLBLM_R_X103Y116_SLICE_X162Y116_A5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_BMUX = CLBLM_R_X103Y116_SLICE_X162Y116_B5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_DMUX = CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A = CLBLM_R_X103Y116_SLICE_X163Y116_AO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B = CLBLM_R_X103Y116_SLICE_X163Y116_BO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C = CLBLM_R_X103Y116_SLICE_X163Y116_CO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D = CLBLM_R_X103Y116_SLICE_X163Y116_DO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_AMUX = CLBLM_R_X103Y116_SLICE_X163Y116_A5Q;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_BMUX = CLBLM_R_X103Y116_SLICE_X163Y116_B5Q;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_CMUX = CLBLM_R_X103Y116_SLICE_X163Y116_CO5;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A = CLBLM_R_X103Y117_SLICE_X162Y117_AO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B = CLBLM_R_X103Y117_SLICE_X162Y117_BO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C = CLBLM_R_X103Y117_SLICE_X162Y117_CO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D = CLBLM_R_X103Y117_SLICE_X162Y117_DO6;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A = CLBLM_R_X103Y117_SLICE_X163Y117_AO6;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B = CLBLM_R_X103Y117_SLICE_X163Y117_BO6;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C = CLBLM_R_X103Y117_SLICE_X163Y117_CO6;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D = CLBLM_R_X103Y117_SLICE_X163Y117_DO6;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_A = CLBLM_R_X103Y118_SLICE_X162Y118_AO6;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_B = CLBLM_R_X103Y118_SLICE_X162Y118_BO6;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_C = CLBLM_R_X103Y118_SLICE_X162Y118_CO6;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_D = CLBLM_R_X103Y118_SLICE_X162Y118_DO6;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_AMUX = CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_BMUX = CLBLM_R_X103Y118_SLICE_X162Y118_B5Q;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_CMUX = CLBLM_R_X103Y118_SLICE_X162Y118_CO5;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_A = CLBLM_R_X103Y118_SLICE_X163Y118_AO6;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_B = CLBLM_R_X103Y118_SLICE_X163Y118_BO6;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_C = CLBLM_R_X103Y118_SLICE_X163Y118_CO6;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_D = CLBLM_R_X103Y118_SLICE_X163Y118_DO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A = CLBLM_R_X103Y119_SLICE_X162Y119_AO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B = CLBLM_R_X103Y119_SLICE_X162Y119_BO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C = CLBLM_R_X103Y119_SLICE_X162Y119_CO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D = CLBLM_R_X103Y119_SLICE_X162Y119_DO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_DMUX = CLBLM_R_X103Y119_SLICE_X162Y119_DO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A = CLBLM_R_X103Y119_SLICE_X163Y119_AO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B = CLBLM_R_X103Y119_SLICE_X163Y119_BO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C = CLBLM_R_X103Y119_SLICE_X163Y119_CO6;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D = CLBLM_R_X103Y119_SLICE_X163Y119_DO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A = CLBLM_R_X103Y122_SLICE_X162Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B = CLBLM_R_X103Y122_SLICE_X162Y122_BO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C = CLBLM_R_X103Y122_SLICE_X162Y122_CO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D = CLBLM_R_X103Y122_SLICE_X162Y122_DO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A = CLBLM_R_X103Y122_SLICE_X163Y122_AO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B = CLBLM_R_X103Y122_SLICE_X163Y122_BO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C = CLBLM_R_X103Y122_SLICE_X163Y122_CO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D = CLBLM_R_X103Y122_SLICE_X163Y122_DO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X102Y107_SLICE_X160Y107_A5Q;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X102Y107_SLICE_X160Y107_AQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X102Y107_SLICE_X160Y107_BQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLM_R_X103Y109_SLICE_X163Y109_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = 1'b0;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = 1'b0;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = 1'b0;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = 1'b0;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = 1'b0;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = 1'b0;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = 1'b0;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = 1'b0;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = 1'b0;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = 1'b0;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = 1'b0;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = 1'b0;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = 1'b0;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = 1'b0;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = 1'b0;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = 1'b0;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = 1'b0;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = 1'b0;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = 1'b0;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = 1'b0;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = 1'b0;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = 1'b0;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = 1'b0;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLM_R_X103Y119_SLICE_X162Y119_BQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = 1'b0;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLM_R_X103Y108_SLICE_X162Y108_CO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = 1'b0;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = 1'b0;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_OQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_TQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_OQ = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_OQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_TQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_OQ = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_OQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_TQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_OQ = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_OQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_TQ = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_OQ = CLBLM_R_X103Y122_SLICE_X163Y122_AQ;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_TQ = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_OQ = 1'b0;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_TQ = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_OQ = 1'b0;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_OQ = 1'b0;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_TQ = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_OQ = 1'b0;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_OQ = 1'b0;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_TQ = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_OQ = 1'b0;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_OQ = 1'b0;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_TQ = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_OQ = 1'b0;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_OQ = CLBLL_L_X102Y107_SLICE_X160Y107_CQ;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_TQ = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_OQ = 1'b0;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_OQ = CLBLM_R_X103Y113_SLICE_X162Y113_DQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_TQ = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_OQ = CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_OQ = CLBLM_R_X103Y118_SLICE_X162Y118_AQ;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_TQ = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_OQ = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_OQ = CLBLM_R_X103Y118_SLICE_X162Y118_BQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_TQ = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_OQ = CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_OQ = CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_OQ = 1'b0;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_OQ = CLBLM_R_X103Y116_SLICE_X163Y116_DQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_OQ = 1'b0;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_TQ = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D2 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = 1'b0;
  assign LIOB33_X0Y147_IOB_X0Y147_O = 1'b0;
  assign RIOB33_SING_X105Y149_IOB_X1Y149_O = CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A3 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A4 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_A6 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B3 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B4 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_B6 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C3 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C4 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_C6 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D3 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D4 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X163Y119_D6 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A1 = CLBLM_R_X103Y118_SLICE_X162Y118_CO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A2 = CLBLM_R_X103Y118_SLICE_X162Y118_BQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A3 = CLBLM_R_X103Y118_SLICE_X162Y118_AQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A4 = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A5 = CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_A6 = CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B1 = CLBLM_R_X103Y118_SLICE_X162Y118_CO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B2 = CLBLM_R_X103Y119_SLICE_X162Y119_BQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B3 = CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B4 = CLBLM_R_X103Y119_SLICE_X162Y119_DO6;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B5 = CLBLM_R_X103Y118_SLICE_X162Y118_BQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_B6 = CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C1 = CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C2 = CLBLM_R_X103Y118_SLICE_X162Y118_AQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C3 = CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C4 = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C5 = CLBLM_R_X103Y119_SLICE_X162Y119_BQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_C6 = CLBLM_R_X103Y118_SLICE_X162Y118_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = 1'b0;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D1 = CLBLM_R_X103Y118_SLICE_X162Y118_AQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D2 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D3 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D4 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D5 = 1'b1;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_D6 = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_D1 = CLBLL_L_X102Y107_SLICE_X160Y107_CQ;
  assign CLBLM_R_X103Y119_SLICE_X162Y119_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = 1'b0;
  assign RIOI3_X105Y139_OLOGIC_X1Y140_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOB33_X105Y145_IOB_X1Y146_O = CLBLM_R_X103Y118_SLICE_X162Y118_AQ;
  assign RIOB33_X105Y145_IOB_X1Y145_O = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign LIOB33_X0Y119_IOB_X0Y120_O = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = 1'b1;
  assign RIOI3_X105Y139_OLOGIC_X1Y139_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y138_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_D1 = 1'b0;
  assign RIOI3_TBYTETERM_X105Y137_OLOGIC_X1Y137_T1 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A1 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A3 = CLBLL_L_X102Y115_SLICE_X160Y115_AQ;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A4 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A5 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_A6 = CLBLL_L_X102Y115_SLICE_X161Y115_CQ;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B1 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B2 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B4 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B5 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_B6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C1 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C2 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C4 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C5 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_C6 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D1 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D2 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D4 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D5 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_D6 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X160Y115_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y117_IOB_X1Y117_O = 1'b1;
  assign RIOB33_X105Y117_IOB_X1Y118_O = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A1 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A2 = CLBLL_L_X102Y115_SLICE_X161Y115_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A3 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A5 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_A6 = CLBLL_L_X102Y115_SLICE_X161Y115_AQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_AX = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B1 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B2 = CLBLL_L_X102Y115_SLICE_X161Y115_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B3 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B5 = CLBLL_L_X102Y115_SLICE_X160Y115_AQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_B6 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C1 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C2 = CLBLL_L_X102Y115_SLICE_X161Y115_CQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C3 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C5 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_C6 = CLBLM_R_X103Y115_SLICE_X162Y115_CQ;
  assign LIOB33_X0Y151_IOB_X0Y151_O = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y152_O = 1'b0;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D1 = CLBLL_L_X102Y115_SLICE_X160Y115_AQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D2 = CLBLL_L_X102Y115_SLICE_X161Y115_CQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D3 = 1'b1;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D4 = CLBLL_L_X102Y115_SLICE_X161Y115_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D5 = CLBLL_L_X102Y115_SLICE_X161Y115_AQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_D6 = CLBLM_R_X103Y116_SLICE_X162Y116_BQ;
  assign CLBLL_L_X102Y115_SLICE_X161Y115_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D2 = 1'b1;
  assign RIOB33_X105Y147_IOB_X1Y148_O = CLBLM_R_X103Y118_SLICE_X162Y118_BQ;
  assign RIOB33_X105Y147_IOB_X1Y147_O = CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  assign LIOB33_X0Y121_IOB_X0Y122_O = 1'b0;
  assign LIOB33_X0Y121_IOB_X0Y121_O = 1'b0;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = 1'b0;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = 1'b0;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y126_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_D1 = 1'b0;
  assign RIOI3_X105Y125_OLOGIC_X1Y125_T1 = 1'b1;
  assign RIOB33_X105Y119_IOB_X1Y120_O = 1'b1;
  assign RIOB33_X105Y119_IOB_X1Y119_O = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_D1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y120_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_D1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_OLOGIC_X1Y119_T1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_A6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_AX = CLBLM_R_X103Y108_SLICE_X162Y108_CO5;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_B6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_C6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_D6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X163Y108_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A1 = CLBLM_R_X103Y108_SLICE_X162Y108_B5Q;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A3 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A4 = CLBLM_R_X103Y109_SLICE_X163Y109_CQ;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A5 = CLBLM_R_X103Y108_SLICE_X162Y108_A5Q;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_A6 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y123_O = 1'b0;
  assign LIOB33_X0Y123_IOB_X0Y124_O = 1'b0;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B5 = CLBLM_R_X103Y108_SLICE_X163Y108_AQ;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_B6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C4 = CLBLM_R_X103Y109_SLICE_X163Y109_AQ;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_C6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D1 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D2 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D3 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D4 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D5 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_D6 = 1'b1;
  assign CLBLM_R_X103Y108_SLICE_X162Y108_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOB33_X0Y105_IOB_X0Y106_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOB33_X0Y105_IOB_X0Y105_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y121_IOB_X1Y122_O = 1'b1;
  assign RIOB33_X105Y121_IOB_X1Y121_O = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = 1'b0;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_D1 = CLBLM_R_X103Y113_SLICE_X162Y113_DQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = 1'b0;
  assign RIOI3_X105Y141_OLOGIC_X1Y142_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_D1 = CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = 1'b0;
  assign RIOI3_X105Y141_OLOGIC_X1Y141_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A1 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_A1 = CLBLM_R_X103Y109_SLICE_X163Y109_B5Q;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_A5 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_A6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A3 = CLBLM_R_X103Y122_SLICE_X163Y122_AQ;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A4 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_B1 = CLBLM_R_X103Y109_SLICE_X163Y109_CQ;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_B2 = CLBLM_R_X103Y109_SLICE_X163Y109_BQ;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_B4 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_B5 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_B6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B2 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_C1 = CLBLL_L_X102Y108_SLICE_X161Y108_B5Q;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_C2 = CLBLL_L_X102Y109_SLICE_X161Y109_AQ;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_C3 = CLBLM_R_X103Y109_SLICE_X162Y109_BQ;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_C5 = CLBLM_R_X103Y109_SLICE_X163Y109_B5Q;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_C6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C1 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_D1 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_D2 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_D3 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_D4 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_D5 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_D6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D1 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X163Y109_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A1 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_A1 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_A2 = CLBLM_R_X103Y108_SLICE_X162Y108_BQ;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_A3 = CLBLL_L_X102Y109_SLICE_X160Y109_BQ;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_A4 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_A6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A5 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_B1 = CLBLL_L_X102Y109_SLICE_X160Y109_B5Q;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_B2 = CLBLM_R_X103Y109_SLICE_X162Y109_A5Q;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_B3 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_B4 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_B6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B5 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_C1 = CLBLM_R_X103Y109_SLICE_X163Y109_AQ;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_C2 = CLBLM_R_X103Y109_SLICE_X162Y109_AQ;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_C4 = CLBLL_L_X102Y109_SLICE_X161Y109_B5Q;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_C5 = CLBLM_R_X103Y109_SLICE_X162Y109_B5Q;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_C6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C2 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_C6 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_D1 = CLBLM_R_X103Y109_SLICE_X162Y109_CO5;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_D2 = CLBLL_L_X102Y110_SLICE_X161Y110_B5Q;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_D3 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_D4 = CLBLM_R_X103Y109_SLICE_X162Y109_A5Q;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_D5 = CLBLM_R_X103Y108_SLICE_X163Y108_AQ;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_D6 = CLBLM_R_X103Y109_SLICE_X163Y109_BQ;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D2 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D3 = 1'b1;
  assign CLBLM_R_X103Y109_SLICE_X162Y109_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D5 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_D6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOB33_X105Y139_IOB_X1Y140_O = CLBLL_L_X102Y107_SLICE_X160Y107_CQ;
  assign RIOB33_X105Y123_IOB_X1Y124_O = 1'b1;
  assign RIOB33_X105Y123_IOB_X1Y123_O = CLBLM_R_X103Y122_SLICE_X163Y122_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = 1'b0;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = 1'b0;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = 1'b0;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = 1'b0;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_D1 = 1'b0;
  assign LIOB33_X0Y127_IOB_X0Y128_O = 1'b0;
  assign LIOB33_X0Y127_IOB_X0Y127_O = 1'b0;
  assign RIOI3_X105Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_A1 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_A2 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_A3 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_A4 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_A5 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_D1 = 1'b0;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_B1 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_B2 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_B3 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_B4 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_B5 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y132_T1 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_C1 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_C2 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_C3 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_C4 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_C5 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_D1 = 1'b0;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_D1 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_D2 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_D3 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_D4 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_D5 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X163Y110_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_OLOGIC_X1Y131_T1 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_A1 = CLBLM_R_X103Y110_SLICE_X162Y110_B5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_A2 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_A3 = CLBLL_L_X102Y108_SLICE_X161Y108_B5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_A5 = CLBLL_L_X102Y108_SLICE_X161Y108_AQ;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_A6 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_B1 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_B3 = CLBLL_L_X102Y108_SLICE_X161Y108_B5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_B4 = CLBLL_L_X102Y110_SLICE_X161Y110_B5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_B5 = CLBLM_R_X103Y110_SLICE_X162Y110_C5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_B6 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_C1 = CLBLM_R_X103Y109_SLICE_X163Y109_CQ;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_C2 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_C3 = CLBLM_R_X103Y109_SLICE_X163Y109_B5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_C4 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_C6 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_D2 = CLBLM_R_X103Y110_SLICE_X162Y110_CQ;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_D3 = CLBLL_L_X102Y109_SLICE_X160Y109_B5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_D4 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_D5 = CLBLM_R_X103Y110_SLICE_X162Y110_D5Q;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_D6 = 1'b1;
  assign CLBLM_R_X103Y110_SLICE_X162Y110_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y125_IOB_X1Y126_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOB33_X105Y125_IOB_X1Y125_O = 1'b0;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOB33_X0Y129_IOB_X0Y130_O = 1'b0;
  assign LIOB33_X0Y129_IOB_X0Y129_O = 1'b0;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = 1'b0;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X102Y107_SLICE_X160Y107_A5Q;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_A6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = 1'b0;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_AX = CLBLM_R_X103Y111_SLICE_X162Y111_A5Q;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_D1 = CLBLM_R_X103Y118_SLICE_X162Y118_AQ;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_B6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X102Y107_SLICE_X160Y107_AQ;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_D1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_BX = CLBLM_R_X103Y108_SLICE_X162Y108_AQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_C6 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y116_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_D1 = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = 1'b0;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_CX = CLBLM_R_X103Y110_SLICE_X162Y110_DQ;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_D6 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_D1 = 1'b1;
  assign RIOI3_X105Y145_OLOGIC_X1Y145_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_DX = CLBLM_R_X103Y110_SLICE_X162Y110_A5Q;
  assign CLBLM_R_X103Y111_SLICE_X163Y111_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A2 = CLBLL_L_X102Y110_SLICE_X161Y110_B5Q;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A4 = CLBLM_R_X103Y110_SLICE_X162Y110_BQ;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_A6 = 1'b1;
  assign RIOI3_X105Y115_OLOGIC_X1Y115_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = 1'b0;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B1 = CLBLM_R_X103Y111_SLICE_X162Y111_B5Q;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B2 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B3 = CLBLM_R_X103Y111_SLICE_X162Y111_AQ;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B4 = CLBLM_R_X103Y108_SLICE_X163Y108_AQ;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_C6 = 1'b1;
  assign RIOB33_X105Y127_IOB_X1Y127_O = 1'b0;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X102Y107_SLICE_X160Y107_A5Q;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X102Y107_SLICE_X160Y107_AQ;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D1 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D2 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D3 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D4 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D5 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_D6 = 1'b1;
  assign CLBLM_R_X103Y111_SLICE_X162Y111_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_A1 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_A3 = CLBLL_L_X102Y107_SLICE_X160Y107_AQ;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_A4 = CLBLM_R_X103Y119_SLICE_X162Y119_CO6;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_A5 = CLBLL_L_X102Y107_SLICE_X160Y107_A5Q;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_A6 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_B1 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_B3 = CLBLL_L_X102Y107_SLICE_X160Y107_AQ;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_B4 = CLBLM_R_X103Y119_SLICE_X162Y119_CO6;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_B5 = CLBLL_L_X102Y107_SLICE_X160Y107_A5Q;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_B6 = CLBLL_L_X102Y107_SLICE_X160Y107_BQ;
  assign LIOB33_X0Y131_IOB_X0Y132_O = 1'b0;
  assign LIOB33_X0Y131_IOB_X0Y131_O = 1'b0;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_C1 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_C2 = CLBLL_L_X102Y107_SLICE_X160Y107_AQ;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_C3 = CLBLL_L_X102Y107_SLICE_X160Y107_BQ;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_C4 = CLBLL_L_X102Y107_SLICE_X160Y107_A5Q;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_C5 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_C6 = CLBLM_R_X103Y119_SLICE_X162Y119_CO6;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_D1 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_D2 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_D3 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_D4 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_D5 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_D6 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X160Y107_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_A1 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_A2 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_A3 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_A4 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_A5 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_A6 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_B1 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_B2 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_B3 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_B4 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_B5 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_B6 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_C1 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_C2 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_C3 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_C4 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A5 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A6 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_C5 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_C6 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_A4 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B4 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_D1 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_D2 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_D3 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_D4 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_D5 = 1'b1;
  assign CLBLL_L_X102Y107_SLICE_X161Y107_D6 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B6 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C4 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C5 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_C6 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D4 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D5 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = 1'b0;
  assign RIOB33_X105Y129_IOB_X1Y129_O = 1'b0;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOB33_X105Y129_IOB_X1Y130_O = 1'b0;
  assign LIOB33_X0Y103_IOB_X0Y104_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X102Y107_SLICE_X160Y107_BQ;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A1 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A2 = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A5 = CLBLL_L_X102Y108_SLICE_X161Y108_B5Q;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B4 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B5 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = 1'b0;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_D1 = 1'b0;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C4 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C5 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_C6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y130_T1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D1 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D2 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D3 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D4 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D5 = 1'b1;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_D6 = 1'b1;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_D1 = 1'b0;
  assign CLBLM_R_X103Y112_SLICE_X162Y112_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y129_OLOGIC_X1Y129_T1 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_D1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_D1 = 1'b0;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y144_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_D1 = CLBLM_R_X103Y116_SLICE_X163Y116_DQ;
  assign RIOI3_TBYTESRC_X105Y143_OLOGIC_X1Y143_T1 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = 1'b0;
  assign LIOB33_X0Y133_IOB_X0Y133_O = 1'b0;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_A1 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_A2 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_A3 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_A4 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_A5 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_A6 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_B1 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_B2 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_B3 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_B4 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_B5 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_B6 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_C1 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_C2 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_C3 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_C4 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_C5 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_C6 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_D1 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_D2 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_D3 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_D4 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_D5 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X160Y108_D6 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_A1 = CLBLL_L_X102Y109_SLICE_X161Y109_DO6;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_A2 = CLBLL_L_X102Y109_SLICE_X161Y109_CO5;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_A4 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_A5 = CLBLM_R_X103Y109_SLICE_X162Y109_DO6;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_A6 = CLBLL_L_X102Y108_SLICE_X161Y108_CO6;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_B1 = CLBLM_R_X103Y109_SLICE_X162Y109_CQ;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_B2 = CLBLL_L_X102Y110_SLICE_X161Y110_B5Q;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_B4 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_B5 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_B6 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_C1 = CLBLM_R_X103Y109_SLICE_X163Y109_CQ;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_C2 = CLBLL_L_X102Y109_SLICE_X161Y109_AO5;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_C3 = CLBLL_L_X102Y108_SLICE_X161Y108_BQ;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_C4 = CLBLM_R_X103Y109_SLICE_X162Y109_CQ;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_C5 = CLBLL_L_X102Y109_SLICE_X161Y109_BQ;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_C6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A1 = CLBLM_R_X103Y113_SLICE_X162Y113_DQ;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A2 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A4 = CLBLM_R_X103Y113_SLICE_X162Y113_BQ;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A5 = CLBLM_R_X103Y113_SLICE_X163Y113_CQ;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_A6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_AX = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_D1 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_D2 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_D3 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_D4 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_D5 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_D6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B1 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B2 = 1'b1;
  assign CLBLL_L_X102Y108_SLICE_X161Y108_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B4 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B5 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_B6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_BX = CLBLM_R_X103Y113_SLICE_X163Y113_AQ;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C1 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C2 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C5 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_C4 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_CX = CLBLM_R_X103Y113_SLICE_X162Y113_DQ;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D1 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D2 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D4 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D5 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X163Y113_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A1 = CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A2 = CLBLL_L_X102Y112_SLICE_X161Y112_CO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A3 = CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A4 = CLBLM_R_X103Y113_SLICE_X162Y113_AQ;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A5 = CLBLM_R_X103Y113_SLICE_X162Y113_A5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_A6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B1 = CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B2 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B3 = CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B4 = CLBLL_L_X102Y112_SLICE_X161Y112_CO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B5 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_B6 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C1 = CLBLM_R_X103Y113_SLICE_X162Y113_AQ;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C2 = CLBLM_R_X103Y113_SLICE_X162Y113_CQ;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C3 = CLBLM_R_X103Y113_SLICE_X163Y113_AO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C4 = CLBLM_R_X103Y113_SLICE_X162Y113_A5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C5 = CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_C6 = CLBLL_L_X102Y112_SLICE_X161Y112_CO6;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D1 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D2 = CLBLM_R_X103Y113_SLICE_X162Y113_CQ;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D3 = 1'b1;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D4 = CLBLM_R_X103Y113_SLICE_X162Y113_A5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D5 = CLBLM_R_X103Y113_SLICE_X162Y113_B5Q;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_D6 = CLBLM_R_X103Y113_SLICE_X162Y113_AQ;
  assign CLBLM_R_X103Y113_SLICE_X162Y113_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = 1'b0;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_D1 = CLBLM_R_X103Y118_SLICE_X162Y118_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = 1'b0;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_D1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X102Y107_SLICE_X160Y107_BQ;
  assign RIOI3_X105Y147_OLOGIC_X1Y148_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y118_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_D1 = CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_D1 = 1'b1;
  assign RIOI3_X105Y147_OLOGIC_X1Y147_T1 = 1'b1;
  assign RIOI3_X105Y117_OLOGIC_X1Y117_T1 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = 1'b0;
  assign LIOB33_X0Y135_IOB_X0Y135_O = 1'b0;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_A2 = CLBLL_L_X102Y110_SLICE_X160Y110_D5Q;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_A3 = CLBLL_L_X102Y109_SLICE_X161Y109_B5Q;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_A4 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_A5 = CLBLL_L_X102Y109_SLICE_X161Y109_CQ;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_A6 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_B1 = CLBLM_R_X103Y112_SLICE_X162Y112_AQ;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_B2 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_B4 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_B5 = CLBLL_L_X102Y108_SLICE_X161Y108_BQ;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_B6 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_C1 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_C2 = CLBLL_L_X102Y109_SLICE_X160Y109_AQ;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_C4 = CLBLL_L_X102Y109_SLICE_X161Y109_CQ;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_C6 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_D1 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_D2 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_D3 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_D4 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_D5 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_D6 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X160Y109_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_A1 = CLBLL_L_X102Y110_SLICE_X161Y110_BQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_A2 = CLBLL_L_X102Y109_SLICE_X160Y109_B5Q;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_A3 = CLBLL_L_X102Y108_SLICE_X161Y108_AQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_A4 = CLBLL_L_X102Y109_SLICE_X161Y109_CQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_A6 = 1'b1;
  assign RIOB33_X105Y133_IOB_X1Y134_O = 1'b0;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_B1 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_B2 = CLBLL_L_X102Y109_SLICE_X160Y109_CQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_B3 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_B5 = CLBLL_L_X102Y108_SLICE_X161Y108_AQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_B6 = 1'b1;
  assign LIOB33_X0Y107_IOB_X0Y107_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLM_R_X103Y108_SLICE_X162Y108_CO6;
  assign RIOB33_X105Y133_IOB_X1Y133_O = 1'b0;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_C1 = CLBLL_L_X102Y108_SLICE_X161Y108_AQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_C2 = CLBLL_L_X102Y109_SLICE_X161Y109_AQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_C3 = CLBLM_R_X103Y109_SLICE_X162Y109_AQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_C4 = CLBLL_L_X102Y110_SLICE_X161Y110_BQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_C6 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_A1 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_A2 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_A3 = CLBLM_R_X103Y114_SLICE_X163Y114_AQ;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_A4 = CLBLM_R_X103Y116_SLICE_X163Y116_B5Q;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_D1 = 1'b1;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_D2 = CLBLM_R_X103Y108_SLICE_X162Y108_BQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_D3 = CLBLM_R_X103Y112_SLICE_X162Y112_AQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_D4 = CLBLL_L_X102Y109_SLICE_X160Y109_CQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_D5 = CLBLM_R_X103Y109_SLICE_X163Y109_CO6;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_D6 = CLBLL_L_X102Y109_SLICE_X160Y109_BQ;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_A6 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_DX = CLBLL_L_X102Y109_SLICE_X160Y109_C5Q;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_B5 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_B6 = CLBLM_R_X103Y115_SLICE_X163Y115_CQ;
  assign CLBLL_L_X102Y109_SLICE_X161Y109_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_B1 = CLBLM_R_X103Y115_SLICE_X163Y115_DQ;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_B2 = CLBLM_R_X103Y115_SLICE_X163Y115_BQ;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_B3 = CLBLM_R_X103Y115_SLICE_X163Y115_AQ;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_B4 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_C1 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_C2 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_C3 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_C4 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_C5 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_C6 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_D1 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_D2 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_D3 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_D4 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_D5 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_D6 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X163Y114_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_A1 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_A2 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_A3 = CLBLM_R_X103Y114_SLICE_X162Y114_AQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_A4 = CLBLM_R_X103Y115_SLICE_X162Y115_AQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_A5 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_A6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_B1 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_B2 = CLBLM_R_X103Y114_SLICE_X162Y114_BQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_B4 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_B5 = CLBLM_R_X103Y114_SLICE_X163Y114_AQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_B6 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_C1 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_C2 = CLBLM_R_X103Y114_SLICE_X162Y114_CQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_C3 = CLBLM_R_X103Y114_SLICE_X162Y114_AQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_C4 = 1'b1;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_C6 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_D1 = CLBLM_R_X103Y114_SLICE_X163Y114_AQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_D2 = CLBLM_R_X103Y114_SLICE_X162Y114_CQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_D3 = CLBLM_R_X103Y114_SLICE_X162Y114_AQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_D4 = CLBLM_R_X103Y114_SLICE_X162Y114_BQ;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_D5 = CLBLM_R_X103Y116_SLICE_X163Y116_B5Q;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_D6 = CLBLL_L_X102Y114_SLICE_X161Y114_AQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X103Y114_SLICE_X162Y114_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOB33_X0Y137_IOB_X0Y138_O = 1'b0;
  assign LIOB33_X0Y137_IOB_X0Y137_O = 1'b0;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = 1'b0;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A5 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = 1'b0;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_A6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_D1 = 1'b0;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = 1'b0;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y134_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B3 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B4 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B5 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_D1 = 1'b0;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_A1 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_A2 = CLBLL_L_X102Y110_SLICE_X160Y110_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_A3 = CLBLL_L_X102Y109_SLICE_X160Y109_BQ;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_A4 = CLBLM_R_X103Y110_SLICE_X162Y110_AQ;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_A6 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_B6 = 1'b1;
  assign RIOI3_X105Y133_OLOGIC_X1Y133_T1 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_B1 = CLBLL_L_X102Y109_SLICE_X161Y109_B5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_B2 = CLBLL_L_X102Y109_SLICE_X160Y109_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_B3 = CLBLL_L_X102Y109_SLICE_X160Y109_BQ;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_B4 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_B6 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_C1 = CLBLL_L_X102Y110_SLICE_X160Y110_C5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_C3 = CLBLL_L_X102Y110_SLICE_X160Y110_BQ;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_C4 = CLBLM_R_X103Y109_SLICE_X162Y109_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_C5 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y126_O = 1'b0;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_X0Y125_IOB_X0Y125_O = 1'b0;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_D2 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_D3 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_D4 = CLBLM_R_X103Y109_SLICE_X162Y109_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_D5 = CLBLL_L_X102Y109_SLICE_X160Y109_B5Q;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_D6 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X160Y110_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_C6 = 1'b1;
  assign RIOB33_X105Y135_IOB_X1Y136_O = 1'b0;
  assign RIOB33_X105Y135_IOB_X1Y135_O = 1'b0;
  assign LIOB33_X0Y109_IOB_X0Y110_O = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLM_R_X103Y109_SLICE_X163Y109_AO5;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_A1 = CLBLL_L_X102Y110_SLICE_X160Y110_DQ;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_A2 = CLBLL_L_X102Y110_SLICE_X161Y110_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_A4 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_A5 = CLBLM_R_X103Y109_SLICE_X163Y109_B5Q;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_A6 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_B2 = CLBLL_L_X102Y109_SLICE_X161Y109_BQ;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_B3 = CLBLM_R_X103Y109_SLICE_X162Y109_B5Q;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_B4 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_B5 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_B6 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_C1 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_C2 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_C3 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_C4 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_C5 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_C6 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_CX = CLBLL_L_X102Y111_SLICE_X161Y111_DQ;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_D1 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_D2 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_D3 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_D4 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_D5 = 1'b1;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_D6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A1 = CLBLM_R_X103Y115_SLICE_X163Y115_CQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A4 = CLBLM_R_X103Y115_SLICE_X163Y115_DQ;
  assign CLBLL_L_X102Y110_SLICE_X161Y110_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A5 = CLBLM_R_X103Y113_SLICE_X163Y113_AO5;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B1 = CLBLM_R_X103Y115_SLICE_X163Y115_CQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B2 = CLBLM_R_X103Y115_SLICE_X163Y115_BQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B3 = CLBLM_R_X103Y115_SLICE_X163Y115_AQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B4 = CLBLM_R_X103Y115_SLICE_X163Y115_DQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B5 = CLBLM_R_X103Y113_SLICE_X163Y113_AO5;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_B6 = CLBLM_R_X103Y116_SLICE_X163Y116_CO6;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D5 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C1 = CLBLM_R_X103Y115_SLICE_X163Y115_BQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C2 = CLBLM_R_X103Y113_SLICE_X163Y113_AO5;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C3 = CLBLM_R_X103Y115_SLICE_X163Y115_DQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C4 = CLBLM_R_X103Y116_SLICE_X163Y116_CO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C5 = CLBLM_R_X103Y115_SLICE_X163Y115_CQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_C6 = CLBLM_R_X103Y115_SLICE_X163Y115_AQ;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_D6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D1 = CLBLM_R_X103Y115_SLICE_X163Y115_BQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D2 = CLBLM_R_X103Y113_SLICE_X163Y113_AO5;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D3 = CLBLM_R_X103Y115_SLICE_X163Y115_DQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D4 = CLBLM_R_X103Y116_SLICE_X163Y116_CO6;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D5 = CLBLM_R_X103Y115_SLICE_X163Y115_CQ;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_D6 = CLBLM_R_X103Y115_SLICE_X163Y115_AQ;
  assign CLBLM_R_X103Y122_SLICE_X163Y122_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A1 = CLBLM_R_X103Y114_SLICE_X162Y114_BQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A2 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A3 = CLBLM_R_X103Y115_SLICE_X162Y115_AQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A5 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_A6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B1 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B2 = CLBLM_R_X103Y115_SLICE_X162Y115_BQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B3 = CLBLL_L_X102Y114_SLICE_X161Y114_AQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B5 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_B6 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C1 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C2 = CLBLM_R_X103Y115_SLICE_X162Y115_CQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C3 = CLBLM_R_X103Y115_SLICE_X162Y115_BQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C4 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C5 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D1 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D2 = CLBLM_R_X103Y115_SLICE_X162Y115_CQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D3 = CLBLM_R_X103Y115_SLICE_X162Y115_AQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D4 = CLBLM_R_X103Y115_SLICE_X162Y115_BQ;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D5 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_D6 = CLBLM_R_X103Y114_SLICE_X162Y114_DO6;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_A6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X162Y115_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B1 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = 1'b0;
  assign LIOB33_X0Y139_IOB_X0Y139_O = 1'b0;
  assign RIOI3_X105Y145_OLOGIC_X1Y146_T1 = 1'b1;
  assign CLBLM_R_X103Y122_SLICE_X162Y122_B6 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A1 = CLBLL_L_X102Y112_SLICE_X160Y112_CQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A2 = CLBLL_L_X102Y111_SLICE_X160Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A3 = CLBLL_L_X102Y111_SLICE_X161Y111_DQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A4 = CLBLL_L_X102Y110_SLICE_X160Y110_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A5 = CLBLL_L_X102Y112_SLICE_X161Y112_AQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_A6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = 1'b0;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_AX = CLBLL_L_X102Y111_SLICE_X160Y111_DQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B1 = CLBLL_L_X102Y112_SLICE_X161Y112_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B2 = CLBLL_L_X102Y111_SLICE_X160Y111_A5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B3 = CLBLL_L_X102Y111_SLICE_X160Y111_DQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B4 = CLBLL_L_X102Y112_SLICE_X160Y112_A5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B5 = CLBLL_L_X102Y111_SLICE_X160Y111_C5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_B6 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_BX = CLBLL_L_X102Y111_SLICE_X160Y111_A5Q;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C1 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C2 = CLBLL_L_X102Y112_SLICE_X160Y112_A5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C3 = CLBLL_L_X102Y112_SLICE_X160Y112_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C4 = CLBLL_L_X102Y110_SLICE_X161Y110_CQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C5 = CLBLL_L_X102Y111_SLICE_X160Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_C6 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOB33_X105Y137_IOB_X1Y138_O = 1'b0;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y137_IOB_X1Y137_O = 1'b0;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = 1'b0;
  assign LIOB33_X0Y111_IOB_X0Y112_O = 1'b0;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_CX = CLBLL_L_X102Y110_SLICE_X161Y110_CQ;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D1 = CLBLL_L_X102Y111_SLICE_X160Y111_AO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D2 = CLBLL_L_X102Y112_SLICE_X160Y112_CO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D3 = CLBLL_L_X102Y112_SLICE_X160Y112_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D4 = CLBLL_L_X102Y111_SLICE_X160Y111_CO6;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D5 = CLBLL_L_X102Y112_SLICE_X160Y112_CQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_D6 = CLBLL_L_X102Y111_SLICE_X160Y111_BO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_DX = CLBLL_L_X102Y111_SLICE_X160Y111_CQ;
  assign CLBLL_L_X102Y111_SLICE_X160Y111_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = 1'b0;
  assign RIOI3_X105Y121_OLOGIC_X1Y122_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_D1 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A1 = CLBLL_L_X102Y111_SLICE_X161Y111_AQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A2 = CLBLL_L_X102Y111_SLICE_X161Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A3 = CLBLL_L_X102Y111_SLICE_X161Y111_CQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A4 = CLBLL_L_X102Y111_SLICE_X160Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A5 = CLBLL_L_X102Y111_SLICE_X160Y111_CQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_A6 = CLBLL_L_X102Y112_SLICE_X160Y112_A5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = 1'b0;
  assign RIOI3_X105Y121_OLOGIC_X1Y121_T1 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_AX = CLBLL_L_X102Y110_SLICE_X160Y110_CQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B1 = CLBLL_L_X102Y111_SLICE_X161Y111_AQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B2 = CLBLL_L_X102Y112_SLICE_X160Y112_A5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B3 = CLBLL_L_X102Y111_SLICE_X161Y111_CQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B4 = CLBLL_L_X102Y111_SLICE_X160Y111_DQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B5 = CLBLM_R_X103Y111_SLICE_X163Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_B6 = CLBLL_L_X102Y111_SLICE_X160Y111_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_BX = CLBLM_R_X103Y111_SLICE_X162Y111_BQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C1 = CLBLL_L_X102Y111_SLICE_X160Y111_AQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C2 = CLBLL_L_X102Y111_SLICE_X160Y111_A5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C3 = CLBLM_R_X103Y111_SLICE_X163Y111_CQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C4 = CLBLL_L_X102Y112_SLICE_X161Y112_AQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C5 = CLBLL_L_X102Y112_SLICE_X161Y112_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_C6 = CLBLM_R_X103Y111_SLICE_X163Y111_AQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_CX = CLBLL_L_X102Y110_SLICE_X161Y110_AQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D1 = 1'b1;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D2 = CLBLM_R_X103Y111_SLICE_X163Y111_DQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D3 = CLBLL_L_X102Y111_SLICE_X160Y111_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D4 = CLBLL_L_X102Y111_SLICE_X161Y111_CO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D5 = CLBLL_L_X102Y109_SLICE_X161Y109_DQ;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_D6 = CLBLL_L_X102Y111_SLICE_X161Y111_DQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A1 = CLBLM_R_X103Y116_SLICE_X163Y116_AQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A2 = CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_DX = CLBLL_L_X102Y112_SLICE_X161Y112_B5Q;
  assign CLBLL_L_X102Y111_SLICE_X161Y111_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A3 = CLBLM_R_X103Y116_SLICE_X163Y116_A5Q;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A4 = CLBLM_R_X103Y117_SLICE_X162Y117_BO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A5 = CLBLM_R_X103Y116_SLICE_X162Y116_CQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_A6 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B1 = CLBLM_R_X103Y116_SLICE_X163Y116_BQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B2 = CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B3 = CLBLM_R_X103Y116_SLICE_X163Y116_AQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B4 = CLBLM_R_X103Y117_SLICE_X162Y117_BO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B5 = CLBLM_R_X103Y116_SLICE_X162Y116_CQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_B6 = CLBLM_R_X103Y116_SLICE_X163Y116_A5Q;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_BX = CLBLM_R_X103Y116_SLICE_X163Y116_CO5;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C1 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C2 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C3 = CLBLM_R_X103Y117_SLICE_X162Y117_CO6;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C5 = CLBLM_R_X103Y116_SLICE_X163Y116_B5Q;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_C6 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D1 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D2 = CLBLM_R_X103Y116_SLICE_X163Y116_BQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D3 = CLBLM_R_X103Y116_SLICE_X163Y116_A5Q;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D4 = CLBLM_R_X103Y116_SLICE_X162Y116_CQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D5 = CLBLM_R_X103Y116_SLICE_X163Y116_AQ;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_D6 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X163Y116_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A1 = CLBLL_L_X102Y115_SLICE_X161Y115_AQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A2 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A3 = CLBLM_R_X103Y116_SLICE_X162Y116_AQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A5 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_A6 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_AX = CLBLM_R_X103Y117_SLICE_X162Y117_BO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B1 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B2 = CLBLM_R_X103Y116_SLICE_X162Y116_BQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B3 = CLBLM_R_X103Y116_SLICE_X162Y116_AQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B5 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_B6 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_BX = CLBLM_R_X103Y116_SLICE_X163Y116_DQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C1 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C2 = CLBLM_R_X103Y116_SLICE_X162Y116_CQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C3 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C4 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C5 = CLBLM_R_X103Y116_SLICE_X162Y116_DO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_C6 = CLBLM_R_X103Y117_SLICE_X162Y117_BO6;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D1 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D2 = 1'b1;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D3 = CLBLM_R_X103Y116_SLICE_X163Y116_DQ;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D4 = CLBLM_R_X103Y116_SLICE_X162Y116_A5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D5 = CLBLM_R_X103Y116_SLICE_X162Y116_B5Q;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_D6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = 1'b0;
  assign LIOB33_X0Y141_IOB_X0Y142_O = 1'b0;
  assign CLBLM_R_X103Y116_SLICE_X162Y116_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y112_SLICE_X163Y112_B5 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLM_R_X103Y119_SLICE_X162Y119_BQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A2 = CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A3 = CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A4 = CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A5 = CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_A6 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign LIOB33_X0Y113_IOB_X0Y114_O = 1'b0;
  assign LIOB33_X0Y113_IOB_X0Y113_O = 1'b0;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_AX = CLBLL_L_X102Y112_SLICE_X161Y112_AQ;
  assign RIOB33_X105Y139_IOB_X1Y139_O = 1'b0;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B2 = CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B3 = CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B4 = CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B5 = CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_B6 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_BX = CLBLL_L_X102Y112_SLICE_X160Y112_CQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C1 = CLBLL_L_X102Y112_SLICE_X160Y112_C5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C2 = CLBLL_L_X102Y111_SLICE_X160Y111_CQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C3 = CLBLL_L_X102Y112_SLICE_X160Y112_DQ;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C4 = CLBLL_L_X102Y111_SLICE_X160Y111_B5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C5 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_C6 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_CX = CLBLL_L_X102Y111_SLICE_X160Y111_C5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D1 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D2 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D3 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D4 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D5 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_D6 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_DX = CLBLL_L_X102Y112_SLICE_X160Y112_C5Q;
  assign CLBLL_L_X102Y112_SLICE_X160Y112_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A1 = CLBLL_L_X102Y111_SLICE_X160Y111_DO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A2 = CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A3 = CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A4 = CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A5 = CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_A6 = CLBLL_L_X102Y112_SLICE_X161Y112_A5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = 1'b0;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_AX = CLBLL_L_X102Y110_SLICE_X160Y110_AQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B2 = CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B3 = CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B4 = CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B5 = CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_B6 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_BX = CLBLL_L_X102Y111_SLICE_X160Y111_B5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C1 = CLBLL_L_X102Y111_SLICE_X161Y111_AO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C2 = CLBLL_L_X102Y111_SLICE_X161Y111_DO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C3 = CLBLL_L_X102Y111_SLICE_X160Y111_DO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C4 = CLBLL_L_X102Y112_SLICE_X161Y112_A5Q;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C5 = CLBLL_L_X102Y112_SLICE_X161Y112_DO6;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_C6 = CLBLL_L_X102Y111_SLICE_X161Y111_BO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = 1'b0;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_D1 = 1'b0;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D1 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D2 = CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D3 = CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D4 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D5 = CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_D6 = CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y135_OLOGIC_X1Y136_T1 = 1'b1;
  assign CLBLL_L_X102Y112_SLICE_X161Y112_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A1 = CLBLM_R_X103Y118_SLICE_X162Y118_B5Q;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A2 = CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A4 = CLBLM_R_X103Y118_SLICE_X163Y118_BQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_A6 = CLBLM_R_X103Y117_SLICE_X163Y117_AQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLM_R_X103Y108_SLICE_X162Y108_CO6;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_D1 = 1'b0;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B1 = CLBLM_R_X103Y118_SLICE_X162Y118_B5Q;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B2 = CLBLM_R_X103Y117_SLICE_X163Y117_BQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B4 = CLBLM_R_X103Y118_SLICE_X163Y118_BQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_B6 = CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  assign RIOI3_X105Y135_OLOGIC_X1Y135_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C2 = CLBLM_R_X103Y117_SLICE_X163Y117_CQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C3 = CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C4 = CLBLM_R_X103Y118_SLICE_X163Y118_BQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C5 = CLBLM_R_X103Y118_SLICE_X162Y118_B5Q;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_C6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D1 = CLBLM_R_X103Y117_SLICE_X162Y117_AQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D2 = CLBLM_R_X103Y117_SLICE_X163Y117_CQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D3 = CLBLM_R_X103Y117_SLICE_X163Y117_BQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D4 = CLBLM_R_X103Y117_SLICE_X163Y117_AQ;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D5 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X163Y117_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A1 = CLBLM_R_X103Y118_SLICE_X162Y118_B5Q;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A3 = CLBLM_R_X103Y117_SLICE_X162Y117_AQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A4 = CLBLM_R_X103Y118_SLICE_X163Y118_BQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_A6 = CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  assign LIOB33_X0Y143_IOB_X0Y143_O = 1'b0;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B1 = CLBLM_R_X103Y115_SLICE_X162Y115_DO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B2 = CLBLM_R_X103Y116_SLICE_X163Y116_CO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B3 = CLBLM_R_X103Y116_SLICE_X162Y116_AQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B4 = CLBLM_R_X103Y116_SLICE_X162Y116_BQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B5 = CLBLM_R_X103Y114_SLICE_X163Y114_BO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_B6 = CLBLL_L_X102Y115_SLICE_X161Y115_DO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C1 = CLBLM_R_X103Y116_SLICE_X162Y116_AQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C2 = CLBLM_R_X103Y115_SLICE_X162Y115_DO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C3 = CLBLL_L_X102Y115_SLICE_X161Y115_DO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C4 = CLBLM_R_X103Y114_SLICE_X163Y114_BO6;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C5 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_C6 = CLBLM_R_X103Y116_SLICE_X162Y116_BQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOB33_X105Y131_IOB_X1Y132_O = 1'b0;
  assign RIOB33_X105Y131_IOB_X1Y131_O = 1'b0;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D1 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D2 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D3 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D4 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D5 = 1'b1;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_D6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLM_R_X103Y119_SLICE_X162Y119_BQ;
  assign CLBLM_R_X103Y117_SLICE_X162Y117_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y141_IOB_X1Y142_O = CLBLM_R_X103Y113_SLICE_X162Y113_DQ;
  assign RIOB33_X105Y141_IOB_X1Y141_O = CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = 1'b0;
  assign LIOB33_X0Y115_IOB_X0Y115_O = 1'b0;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = 1'b0;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A5 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_A6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B5 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_B6 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C5 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_C6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = 1'b0;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D5 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X160Y113_D6 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A1 = CLBLL_L_X102Y113_SLICE_X161Y113_AQ;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A3 = CLBLL_L_X102Y112_SLICE_X161Y112_BQ;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A4 = CLBLL_L_X102Y112_SLICE_X160Y112_BQ;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A5 = CLBLL_L_X102Y112_SLICE_X160Y112_AQ;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_A6 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B5 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_B6 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C5 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_C6 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D1 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D2 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D3 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D4 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D5 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_D6 = 1'b1;
  assign CLBLL_L_X102Y113_SLICE_X161Y113_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_A1 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_A2 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_A3 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_A4 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_A5 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_A6 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_AX = CLBLM_R_X103Y118_SLICE_X162Y118_CO5;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_B1 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_B2 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_B3 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_B4 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_B5 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_B6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = 1'b0;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_BX = CLBLM_R_X103Y118_SLICE_X163Y118_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_C1 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_C2 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_C3 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_C4 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_C5 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_C6 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y145_O = 1'b0;
  assign LIOB33_X0Y145_IOB_X0Y146_O = 1'b0;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = 1'b0;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_D1 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_D2 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_D3 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_D4 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_D5 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_D6 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X163Y118_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLM_R_X103Y109_SLICE_X163Y109_AO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_D1 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_A1 = CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_A2 = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_A3 = CLBLM_R_X103Y118_SLICE_X162Y118_AQ;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_A4 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_A6 = 1'b1;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = 1'b0;
  assign RIOI3_X105Y123_OLOGIC_X1Y124_T1 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_B1 = CLBLM_R_X103Y118_SLICE_X162Y118_BQ;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_B2 = CLBLM_R_X103Y112_SLICE_X162Y112_A5Q;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_B3 = CLBLM_R_X103Y118_SLICE_X162Y118_AQ;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_B4 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_B6 = CLBLM_R_X103Y118_SLICE_X162Y118_A5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_D1 = CLBLM_R_X103Y122_SLICE_X163Y122_AQ;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_BX = CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_C2 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_C3 = CLBLM_R_X103Y117_SLICE_X163Y117_DQ;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_C4 = CLBLL_L_X102Y115_SLICE_X161Y115_A5Q;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_C5 = CLBLM_R_X103Y118_SLICE_X162Y118_B5Q;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_C6 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A2 = CLBLM_R_X103Y115_SLICE_X163Y115_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = 1'b0;
  assign RIOI3_X105Y123_OLOGIC_X1Y123_T1 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A3 = CLBLM_R_X103Y115_SLICE_X163Y115_AQ;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_D1 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_D2 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_D3 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_D4 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_D5 = 1'b1;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X103Y115_SLICE_X163Y115_A6 = CLBLM_R_X103Y116_SLICE_X163Y116_CO6;
  assign CLBLM_R_X103Y118_SLICE_X162Y118_SR = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y143_IOB_X1Y144_O = 1'b0;
  assign RIOB33_X105Y143_IOB_X1Y143_O = CLBLM_R_X103Y116_SLICE_X163Y116_DQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOB33_X0Y117_IOB_X0Y117_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A2 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_A6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B2 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_B6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C2 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_C6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D2 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X160Y114_D6 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign RIOB33_X105Y115_IOB_X1Y116_O = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A2 = CLBLM_R_X103Y114_SLICE_X162Y114_CQ;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A3 = CLBLL_L_X102Y114_SLICE_X161Y114_AQ;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A4 = CLBLM_R_X103Y113_SLICE_X163Y113_BQ;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_A6 = CLBLM_R_X103Y115_SLICE_X162Y115_A5Q;
  assign RIOB33_X105Y115_IOB_X1Y115_O = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_D1 = CLBLM_R_X103Y119_SLICE_X162Y119_AQ;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B2 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_B6 = 1'b1;
  assign RIOI3_SING_X105Y149_OLOGIC_X1Y149_T1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C1 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C2 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C3 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C4 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C5 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_C6 = 1'b1;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X102Y114_SLICE_X161Y114_D1 = 1'b1;
endmodule
