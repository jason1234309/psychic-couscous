module top(
  input LIOB33_SING_X0Y150_IOB_X0Y150_IPAD,
  input LIOB33_SING_X0Y199_IOB_X0Y199_IPAD,
  input LIOB33_SING_X0Y200_IOB_X0Y200_IPAD,
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y151_IOB_X0Y151_IPAD,
  input LIOB33_X0Y151_IOB_X0Y152_IPAD,
  input LIOB33_X0Y153_IOB_X0Y153_IPAD,
  input LIOB33_X0Y153_IOB_X0Y154_IPAD,
  input LIOB33_X0Y155_IOB_X0Y155_IPAD,
  input LIOB33_X0Y155_IOB_X0Y156_IPAD,
  input LIOB33_X0Y157_IOB_X0Y157_IPAD,
  input LIOB33_X0Y157_IOB_X0Y158_IPAD,
  input LIOB33_X0Y159_IOB_X0Y159_IPAD,
  input LIOB33_X0Y159_IOB_X0Y160_IPAD,
  input LIOB33_X0Y161_IOB_X0Y161_IPAD,
  input LIOB33_X0Y161_IOB_X0Y162_IPAD,
  input LIOB33_X0Y163_IOB_X0Y163_IPAD,
  input LIOB33_X0Y163_IOB_X0Y164_IPAD,
  input LIOB33_X0Y165_IOB_X0Y165_IPAD,
  input LIOB33_X0Y165_IOB_X0Y166_IPAD,
  input LIOB33_X0Y167_IOB_X0Y167_IPAD,
  input LIOB33_X0Y167_IOB_X0Y168_IPAD,
  input LIOB33_X0Y169_IOB_X0Y169_IPAD,
  input LIOB33_X0Y169_IOB_X0Y170_IPAD,
  input LIOB33_X0Y171_IOB_X0Y171_IPAD,
  input LIOB33_X0Y171_IOB_X0Y172_IPAD,
  input LIOB33_X0Y173_IOB_X0Y173_IPAD,
  input LIOB33_X0Y173_IOB_X0Y174_IPAD,
  input LIOB33_X0Y175_IOB_X0Y175_IPAD,
  input LIOB33_X0Y175_IOB_X0Y176_IPAD,
  input LIOB33_X0Y177_IOB_X0Y177_IPAD,
  input LIOB33_X0Y177_IOB_X0Y178_IPAD,
  input LIOB33_X0Y179_IOB_X0Y179_IPAD,
  input LIOB33_X0Y179_IOB_X0Y180_IPAD,
  input LIOB33_X0Y181_IOB_X0Y181_IPAD,
  input LIOB33_X0Y181_IOB_X0Y182_IPAD,
  input LIOB33_X0Y183_IOB_X0Y183_IPAD,
  input LIOB33_X0Y183_IOB_X0Y184_IPAD,
  input LIOB33_X0Y185_IOB_X0Y185_IPAD,
  input LIOB33_X0Y185_IOB_X0Y186_IPAD,
  input LIOB33_X0Y187_IOB_X0Y187_IPAD,
  input LIOB33_X0Y187_IOB_X0Y188_IPAD,
  input LIOB33_X0Y189_IOB_X0Y189_IPAD,
  input LIOB33_X0Y189_IOB_X0Y190_IPAD,
  input LIOB33_X0Y191_IOB_X0Y191_IPAD,
  input LIOB33_X0Y191_IOB_X0Y192_IPAD,
  input LIOB33_X0Y193_IOB_X0Y193_IPAD,
  input LIOB33_X0Y193_IOB_X0Y194_IPAD,
  input LIOB33_X0Y195_IOB_X0Y195_IPAD,
  input LIOB33_X0Y195_IOB_X0Y196_IPAD,
  input LIOB33_X0Y197_IOB_X0Y197_IPAD,
  input LIOB33_X0Y197_IOB_X0Y198_IPAD,
  input LIOB33_X0Y201_IOB_X0Y201_IPAD,
  input LIOB33_X0Y201_IOB_X0Y202_IPAD,
  input LIOB33_X0Y203_IOB_X0Y203_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input LIOB33_X0Y79_IOB_X0Y80_IPAD,
  input LIOB33_X0Y81_IOB_X0Y81_IPAD,
  input LIOB33_X0Y81_IOB_X0Y82_IPAD,
  input LIOB33_X0Y83_IOB_X0Y83_IPAD,
  input LIOB33_X0Y83_IOB_X0Y84_IPAD,
  input LIOB33_X0Y85_IOB_X0Y85_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_SING_X105Y150_IOB_X1Y150_IPAD,
  input RIOB33_SING_X105Y199_IOB_X1Y199_IPAD,
  input RIOB33_SING_X105Y50_IOB_X1Y50_IPAD,
  input RIOB33_SING_X105Y99_IOB_X1Y99_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  input RIOB33_X105Y151_IOB_X1Y151_IPAD,
  input RIOB33_X105Y151_IOB_X1Y152_IPAD,
  input RIOB33_X105Y153_IOB_X1Y153_IPAD,
  input RIOB33_X105Y153_IOB_X1Y154_IPAD,
  input RIOB33_X105Y155_IOB_X1Y155_IPAD,
  input RIOB33_X105Y155_IOB_X1Y156_IPAD,
  input RIOB33_X105Y157_IOB_X1Y157_IPAD,
  input RIOB33_X105Y157_IOB_X1Y158_IPAD,
  input RIOB33_X105Y159_IOB_X1Y159_IPAD,
  input RIOB33_X105Y159_IOB_X1Y160_IPAD,
  input RIOB33_X105Y161_IOB_X1Y161_IPAD,
  input RIOB33_X105Y161_IOB_X1Y162_IPAD,
  input RIOB33_X105Y163_IOB_X1Y163_IPAD,
  input RIOB33_X105Y163_IOB_X1Y164_IPAD,
  input RIOB33_X105Y165_IOB_X1Y165_IPAD,
  input RIOB33_X105Y165_IOB_X1Y166_IPAD,
  input RIOB33_X105Y167_IOB_X1Y167_IPAD,
  input RIOB33_X105Y167_IOB_X1Y168_IPAD,
  input RIOB33_X105Y169_IOB_X1Y169_IPAD,
  input RIOB33_X105Y169_IOB_X1Y170_IPAD,
  input RIOB33_X105Y171_IOB_X1Y171_IPAD,
  input RIOB33_X105Y171_IOB_X1Y172_IPAD,
  input RIOB33_X105Y173_IOB_X1Y173_IPAD,
  input RIOB33_X105Y173_IOB_X1Y174_IPAD,
  input RIOB33_X105Y175_IOB_X1Y175_IPAD,
  input RIOB33_X105Y175_IOB_X1Y176_IPAD,
  input RIOB33_X105Y177_IOB_X1Y177_IPAD,
  input RIOB33_X105Y177_IOB_X1Y178_IPAD,
  input RIOB33_X105Y179_IOB_X1Y179_IPAD,
  input RIOB33_X105Y179_IOB_X1Y180_IPAD,
  input RIOB33_X105Y181_IOB_X1Y181_IPAD,
  input RIOB33_X105Y181_IOB_X1Y182_IPAD,
  input RIOB33_X105Y183_IOB_X1Y183_IPAD,
  input RIOB33_X105Y183_IOB_X1Y184_IPAD,
  input RIOB33_X105Y185_IOB_X1Y185_IPAD,
  input RIOB33_X105Y185_IOB_X1Y186_IPAD,
  input RIOB33_X105Y187_IOB_X1Y187_IPAD,
  input RIOB33_X105Y187_IOB_X1Y188_IPAD,
  input RIOB33_X105Y189_IOB_X1Y189_IPAD,
  input RIOB33_X105Y189_IOB_X1Y190_IPAD,
  input RIOB33_X105Y191_IOB_X1Y191_IPAD,
  input RIOB33_X105Y191_IOB_X1Y192_IPAD,
  input RIOB33_X105Y193_IOB_X1Y193_IPAD,
  input RIOB33_X105Y193_IOB_X1Y194_IPAD,
  input RIOB33_X105Y195_IOB_X1Y195_IPAD,
  input RIOB33_X105Y195_IOB_X1Y196_IPAD,
  input RIOB33_X105Y197_IOB_X1Y197_IPAD,
  input RIOB33_X105Y197_IOB_X1Y198_IPAD,
  input RIOB33_X105Y51_IOB_X1Y51_IPAD,
  input RIOB33_X105Y51_IOB_X1Y52_IPAD,
  input RIOB33_X105Y53_IOB_X1Y53_IPAD,
  input RIOB33_X105Y53_IOB_X1Y54_IPAD,
  input RIOB33_X105Y55_IOB_X1Y55_IPAD,
  input RIOB33_X105Y55_IOB_X1Y56_IPAD,
  input RIOB33_X105Y57_IOB_X1Y57_IPAD,
  input RIOB33_X105Y57_IOB_X1Y58_IPAD,
  input RIOB33_X105Y59_IOB_X1Y59_IPAD,
  input RIOB33_X105Y59_IOB_X1Y60_IPAD,
  input RIOB33_X105Y61_IOB_X1Y61_IPAD,
  input RIOB33_X105Y61_IOB_X1Y62_IPAD,
  input RIOB33_X105Y63_IOB_X1Y63_IPAD,
  input RIOB33_X105Y63_IOB_X1Y64_IPAD,
  input RIOB33_X105Y65_IOB_X1Y65_IPAD,
  input RIOB33_X105Y65_IOB_X1Y66_IPAD,
  input RIOB33_X105Y67_IOB_X1Y67_IPAD,
  input RIOB33_X105Y67_IOB_X1Y68_IPAD,
  input RIOB33_X105Y69_IOB_X1Y69_IPAD,
  input RIOB33_X105Y69_IOB_X1Y70_IPAD,
  input RIOB33_X105Y71_IOB_X1Y71_IPAD,
  input RIOB33_X105Y71_IOB_X1Y72_IPAD,
  input RIOB33_X105Y73_IOB_X1Y73_IPAD,
  input RIOB33_X105Y73_IOB_X1Y74_IPAD,
  input RIOB33_X105Y75_IOB_X1Y75_IPAD,
  input RIOB33_X105Y75_IOB_X1Y76_IPAD,
  input RIOB33_X105Y77_IOB_X1Y77_IPAD,
  input RIOB33_X105Y77_IOB_X1Y78_IPAD,
  input RIOB33_X105Y79_IOB_X1Y79_IPAD,
  input RIOB33_X105Y79_IOB_X1Y80_IPAD,
  input RIOB33_X105Y81_IOB_X1Y81_IPAD,
  input RIOB33_X105Y81_IOB_X1Y82_IPAD,
  input RIOB33_X105Y83_IOB_X1Y83_IPAD,
  input RIOB33_X105Y83_IOB_X1Y84_IPAD,
  input RIOB33_X105Y85_IOB_X1Y85_IPAD,
  input RIOB33_X105Y85_IOB_X1Y86_IPAD,
  input RIOB33_X105Y87_IOB_X1Y87_IPAD,
  input RIOB33_X105Y87_IOB_X1Y88_IPAD,
  input RIOB33_X105Y89_IOB_X1Y89_IPAD,
  input RIOB33_X105Y89_IOB_X1Y90_IPAD,
  input RIOB33_X105Y91_IOB_X1Y91_IPAD,
  input RIOB33_X105Y91_IOB_X1Y92_IPAD,
  input RIOB33_X105Y93_IOB_X1Y93_IPAD,
  input RIOB33_X105Y93_IOB_X1Y94_IPAD,
  input RIOB33_X105Y95_IOB_X1Y95_IPAD,
  input RIOB33_X105Y95_IOB_X1Y96_IPAD,
  input RIOB33_X105Y97_IOB_X1Y97_IPAD,
  input RIOB33_X105Y97_IOB_X1Y98_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y99_IOB_X0Y99_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y85_IOB_X0Y86_OPAD,
  output LIOB33_X0Y87_IOB_X0Y87_OPAD,
  output LIOB33_X0Y87_IOB_X0Y88_OPAD,
  output LIOB33_X0Y89_IOB_X0Y89_OPAD,
  output LIOB33_X0Y89_IOB_X0Y90_OPAD,
  output LIOB33_X0Y91_IOB_X0Y91_OPAD,
  output LIOB33_X0Y91_IOB_X0Y92_OPAD,
  output LIOB33_X0Y93_IOB_X0Y93_OPAD,
  output LIOB33_X0Y93_IOB_X0Y94_OPAD,
  output LIOB33_X0Y95_IOB_X0Y95_OPAD,
  output LIOB33_X0Y95_IOB_X0Y96_OPAD,
  output LIOB33_X0Y97_IOB_X0Y97_OPAD,
  output LIOB33_X0Y97_IOB_X0Y98_OPAD
  );
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BMUX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CLK;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CLK;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CLK;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BQ;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CLK;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BQ;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CLK;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AQ;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BQ;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BX;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CLK;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CLK;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AQ;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_AX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BQ;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_BX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CLK;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CQ;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_CX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DQ;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_DX;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X0Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_A_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_B_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_C_XOR;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D1;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D2;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D3;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D4;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO5;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_CY;
  wire [0:0] CLBLL_L_X2Y123_SLICE_X1Y123_D_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AQ;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_AX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_A_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_BO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_BO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_BQ;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_BX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_B_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_CLK;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_CO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_CQ;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_CX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_C_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_DMUX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_DO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_DQ;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_DX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X0Y124_D_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_AO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_AX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_A_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_BO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_BO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_BQ;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_BX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_B_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_CLK;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_CO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_CQ;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_C_XOR;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D1;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D2;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D3;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D4;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_DO5;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_DQ;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_DX;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D_CY;
  wire [0:0] CLBLL_L_X2Y124_SLICE_X1Y124_D_XOR;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_A;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_A1;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_A2;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_A3;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_A4;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_A5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_A6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_AO5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_AO6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_AX;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_A_CY;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_A_XOR;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_B;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_B1;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_B2;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_B3;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_B4;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_B5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_B6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_BMUX;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_BO5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_BO6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_BX;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_B_CY;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_B_XOR;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_C;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_C1;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_C2;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_C3;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_C4;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_C5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_C6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_CO5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_CO6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_CX;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_C_CY;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_C_XOR;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_D;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_D1;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_D2;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_D3;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_D4;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_D5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_D6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_DO5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_DO6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_D_CY;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_D_XOR;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_F7AMUX_O;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_F7BMUX_O;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X106Y116_F8MUX_O;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_A;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_A1;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_A2;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_A3;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_A4;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_A5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_A6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_AO5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_AO6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_A_CY;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_A_XOR;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_B;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_B1;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_B2;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_B3;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_B4;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_B5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_B6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_BO5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_BO6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_B_CY;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_B_XOR;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_C;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_C1;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_C2;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_C3;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_C4;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_C5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_C6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_CO5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_CO6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_C_CY;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_C_XOR;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_D;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_D1;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_D2;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_D3;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_D4;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_D5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_D6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_DO5;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_DO6;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_D_CY;
  wire [0:0] CLBLL_R_X71Y116_SLICE_X107Y116_D_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_AMUX;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_AO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_AO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_AX;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_A_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_BO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_BO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_B_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_CMUX;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_CO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_CO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_CX;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_C_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_DO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_DO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_D_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_F7AMUX_O;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X106Y117_F7BMUX_O;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_AO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_AO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_A_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_BO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_BO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_B_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_CO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_CO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_C_XOR;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D1;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D2;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D3;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D4;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_DO5;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_DO6;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D_CY;
  wire [0:0] CLBLL_R_X71Y117_SLICE_X107Y117_D_XOR;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_A;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_A1;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_A2;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_A3;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_A4;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_A5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_A6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_AO5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_AO6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_A_CY;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_A_XOR;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_B;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_B1;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_B2;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_B3;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_B4;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_B5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_B6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_BO5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_BO6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_B_CY;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_B_XOR;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_C;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_C1;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_C2;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_C3;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_C4;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_C5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_C6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_CO5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_CO6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_C_CY;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_C_XOR;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_D;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_D1;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_D2;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_D3;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_D4;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_D5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_D6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_DO5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_DO6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_D_CY;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X106Y118_D_XOR;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_A;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_A1;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_A2;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_A3;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_A4;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_A5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_A6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_AO5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_AO6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_AX;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_A_CY;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_A_XOR;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_B;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_B1;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_B2;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_B3;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_B4;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_B5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_B6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_BMUX;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_BO5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_BO6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_BX;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_B_CY;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_B_XOR;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_C;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_C1;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_C2;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_C3;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_C4;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_C5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_C6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_CO5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_CO6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_CX;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_C_CY;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_C_XOR;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_D;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_D1;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_D2;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_D3;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_D4;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_D5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_D6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_DO5;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_DO6;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_D_CY;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_D_XOR;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_F7AMUX_O;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_F7BMUX_O;
  wire [0:0] CLBLL_R_X71Y118_SLICE_X107Y118_F8MUX_O;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_AO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_AO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_A_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_BO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_BO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_B_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_CLK;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_CO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_CO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_C_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_DO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_DO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X106Y119_D_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_AMUX;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_AO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_AO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_AX;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_A_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_BO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_BO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_B_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_CMUX;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_CO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_CO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_CX;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_C_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D1;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D2;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D3;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D4;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_DO5;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_DO6;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D_CY;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_D_XOR;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_F7AMUX_O;
  wire [0:0] CLBLL_R_X71Y119_SLICE_X107Y119_F7BMUX_O;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_A;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_A1;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_A2;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_A3;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_A4;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_A5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_A6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_AMUX;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_AO5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_AO6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_AX;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_A_CY;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_A_XOR;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_B;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_B1;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_B2;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_B3;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_B4;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_B5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_B6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_BO5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_BO6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_B_CY;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_B_XOR;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_C;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_C1;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_C2;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_C3;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_C4;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_C5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_C6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_CMUX;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_CO5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_CO6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_CX;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_C_CY;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_C_XOR;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_D;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_D1;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_D2;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_D3;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_D4;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_D5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_D6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_DO5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_DO6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_D_CY;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_D_XOR;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_F7AMUX_O;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X106Y120_F7BMUX_O;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_A;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_A1;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_A2;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_A3;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_A4;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_A5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_A6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_AO5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_AO6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_A_CY;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_A_XOR;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_B;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_B1;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_B2;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_B3;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_B4;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_B5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_B6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_BO5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_BO6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_B_CY;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_B_XOR;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_C;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_C1;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_C2;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_C3;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_C4;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_C5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_C6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_CO5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_CO6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_C_CY;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_C_XOR;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_D;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_D1;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_D2;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_D3;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_D4;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_D5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_D6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_DO5;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_DO6;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_D_CY;
  wire [0:0] CLBLL_R_X71Y120_SLICE_X107Y120_D_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_AMUX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_AO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_AO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_AX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_A_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_BO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_BO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_B_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_CMUX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_CO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_CO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_CX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_C_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_DO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_DO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_D_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_F7AMUX_O;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X106Y121_F7BMUX_O;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_AO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_AO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_AX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_A_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_BMUX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_BO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_BO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_BX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_B_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_CO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_CO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_CX;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_C_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D1;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D2;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D3;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D4;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_DO5;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_DO6;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D_CY;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_D_XOR;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_F7AMUX_O;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_F7BMUX_O;
  wire [0:0] CLBLL_R_X71Y121_SLICE_X107Y121_F8MUX_O;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_A;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_A1;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_A2;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_A3;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_A4;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_A5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_A6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_AMUX;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_AO5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_AO6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_A_CY;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_A_XOR;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_B;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_B1;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_B2;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_B3;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_B4;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_B5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_B6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_BO5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_BO6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_B_CY;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_B_XOR;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_C;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_C1;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_C2;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_C3;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_C4;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_C5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_C6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_CO5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_CO6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_C_CY;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_C_XOR;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_D;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_D1;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_D2;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_D3;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_D4;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_D5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_D6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_DO5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_DO6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_D_CY;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X106Y122_D_XOR;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_A;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_A1;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_A2;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_A3;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_A4;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_A5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_A6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_AO5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_AO6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_A_CY;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_A_XOR;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_B;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_B1;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_B2;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_B3;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_B4;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_B5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_B6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_BO5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_BO6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_B_CY;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_B_XOR;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_C;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_C1;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_C2;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_C3;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_C4;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_C5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_C6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_CO5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_CO6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_C_CY;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_C_XOR;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_D;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_D1;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_D2;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_D3;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_D4;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_D5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_D6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_DO5;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_DO6;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_D_CY;
  wire [0:0] CLBLL_R_X71Y122_SLICE_X107Y122_D_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_AO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_AO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_A_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_BO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_BO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_B_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_CO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_CO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_C_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_DO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_DO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X106Y125_D_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_AMUX;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_AO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_AO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_AX;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_A_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_BO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_B_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_CO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_C_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D1;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D2;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D3;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D4;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_DO5;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_DO6;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D_CY;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_D_XOR;
  wire [0:0] CLBLL_R_X71Y125_SLICE_X107Y125_F7AMUX_O;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_AO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_AO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_A_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_BO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_BO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_B_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_CO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_C_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_DO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_DO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X106Y126_D_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_AMUX;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_AO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_AO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_AX;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_A_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_BO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_BO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_B_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_CO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_CO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_C_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D1;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D2;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D3;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D4;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_DO5;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_DO6;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D_CY;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_D_XOR;
  wire [0:0] CLBLL_R_X71Y126_SLICE_X107Y126_F7AMUX_O;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_AO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_AO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_A_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_BO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_BO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_B_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_CO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_CO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_C_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_DO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_DO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X106Y127_D_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_AO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_AO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_A_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_BO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_BO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_B_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_CO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_CO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_C_XOR;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D1;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D2;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D3;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D4;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_DO5;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_DO6;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D_CY;
  wire [0:0] CLBLL_R_X71Y127_SLICE_X107Y127_D_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_AMUX;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_AO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_AO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_AQ;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_AX;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_A_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_BO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_BO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_BQ;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_BX;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_B_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_CLK;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_CMUX;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_CO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_C_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_DO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_DO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X106Y128_D_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_AO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_AO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_A_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_BO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_BO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_B_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_CO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_CO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_C_XOR;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D1;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D2;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D3;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D4;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_DO5;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_DO6;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D_CY;
  wire [0:0] CLBLL_R_X71Y128_SLICE_X107Y128_D_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_AO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_AO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_A_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_BO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_BO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_B_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_CO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_CO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_C_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_DO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_DO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X106Y129_D_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_AO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_AO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_A_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_BO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_BO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_B_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_CO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_CO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_C_XOR;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D1;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D2;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D3;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D4;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_DO5;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_DO6;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D_CY;
  wire [0:0] CLBLL_R_X71Y129_SLICE_X107Y129_D_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_AO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_AO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_AX;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_A_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_BO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_BO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_BQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_BX;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_B_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_CLK;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_CO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_CO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_C_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_DO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_DO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X106Y131_D_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AMUX;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_AX;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_A_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_BO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_BO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_BQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_B_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CLK;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CMUX;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CQ;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_CX;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_C_XOR;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D1;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D2;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D3;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D4;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_DO5;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D_CY;
  wire [0:0] CLBLL_R_X71Y131_SLICE_X107Y131_D_XOR;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_A;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_A1;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_A2;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_A3;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_A4;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_A5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_A6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_AO5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_AO6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_AX;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_A_CY;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_A_XOR;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_B;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_B1;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_B2;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_B3;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_B4;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_B5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_B6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_BMUX;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_BO5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_BO6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_BX;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_B_CY;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_B_XOR;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_C;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_C1;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_C2;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_C3;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_C4;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_C5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_C6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_CO5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_CO6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_CX;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_C_CY;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_C_XOR;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_D;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_D1;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_D2;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_D3;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_D4;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_D5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_D6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_DO5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_DO6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_D_CY;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_D_XOR;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X110Y114_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_A;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_A1;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_A2;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_A3;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_A4;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_A5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_A6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_AO5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_AO6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_A_CY;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_A_XOR;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_B;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_B1;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_B2;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_B3;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_B4;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_B5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_B6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_BO5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_BO6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_B_CY;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_B_XOR;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_C;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_C1;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_C2;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_C3;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_C4;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_C5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_C6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_CO5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_CO6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_C_CY;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_C_XOR;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_D;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_D1;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_D2;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_D3;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_D4;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_D5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_D6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_DO5;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_DO6;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_D_CY;
  wire [0:0] CLBLL_R_X73Y114_SLICE_X111Y114_D_XOR;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_A;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_A1;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_A2;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_A3;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_A4;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_A5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_A6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_AMUX;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_AO5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_AO6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_AX;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_A_CY;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_A_XOR;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_B;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_B1;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_B2;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_B3;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_B4;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_B5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_B6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_BO5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_BO6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_B_CY;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_B_XOR;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_C;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_C1;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_C2;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_C3;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_C4;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_C5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_C6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_CO5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_CO6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_C_CY;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_C_XOR;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_D;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_D1;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_D2;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_D3;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_D4;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_D5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_D6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_DO5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_DO6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_D_CY;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_D_XOR;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X110Y115_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_A;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_A1;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_A2;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_A3;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_A4;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_A5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_A6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_AO5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_AO6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_AX;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_A_CY;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_A_XOR;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_B;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_B1;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_B2;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_B3;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_B4;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_B5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_B6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_BMUX;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_BO5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_BO6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_BX;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_B_CY;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_B_XOR;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_C;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_C1;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_C2;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_C3;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_C4;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_C5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_C6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_CO5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_CO6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_CX;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_C_CY;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_C_XOR;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_D;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_D1;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_D2;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_D3;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_D4;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_D5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_D6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_DO5;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_DO6;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_D_CY;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_D_XOR;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y115_SLICE_X111Y115_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_A;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_A1;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_A2;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_A3;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_A4;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_A5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_A6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_AMUX;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_AO5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_AO6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_AX;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_A_CY;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_A_XOR;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_B;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_B1;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_B2;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_B3;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_B4;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_B5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_B6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_BO5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_BO6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_B_CY;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_B_XOR;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_C;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_C1;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_C2;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_C3;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_C4;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_C5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_C6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_CO5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_CO6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_C_CY;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_C_XOR;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_D;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_D1;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_D2;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_D3;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_D4;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_D5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_D6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_DO5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_DO6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_D_CY;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_D_XOR;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X110Y116_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_A;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_A1;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_A2;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_A3;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_A4;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_A5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_A6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_AO5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_AO6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_AX;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_A_CY;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_A_XOR;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_B;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_B1;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_B2;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_B3;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_B4;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_B5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_B6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_BMUX;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_BO5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_BO6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_BX;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_B_CY;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_B_XOR;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_C;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_C1;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_C2;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_C3;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_C4;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_C5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_C6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_CO5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_CO6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_CX;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_C_CY;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_C_XOR;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_D;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_D1;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_D2;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_D3;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_D4;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_D5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_D6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_DO5;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_DO6;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_D_CY;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_D_XOR;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y116_SLICE_X111Y116_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_AO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_AO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_AX;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_A_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_BMUX;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_BO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_BO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_BX;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_B_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_CO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_CO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_CX;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_C_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_DO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_DO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_D_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X110Y118_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_AMUX;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_AO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_AO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_AX;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_A_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_BO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_BO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_B_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_CO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_CO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_C_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D1;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D2;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D3;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D4;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_DO5;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_DO6;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D_CY;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_D_XOR;
  wire [0:0] CLBLL_R_X73Y118_SLICE_X111Y118_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_AO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_AO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_AX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_A_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_BMUX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_BO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_BO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_BX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_B_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_CO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_CX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_C_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_DO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_DO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_D_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X110Y119_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_AMUX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_AO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_AO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_AX;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_A_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_BO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_BO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_B_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_CO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_CO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_C_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D1;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D2;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D3;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D4;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_DO5;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D_CY;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_D_XOR;
  wire [0:0] CLBLL_R_X73Y119_SLICE_X111Y119_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_A;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_A1;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_A2;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_A3;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_A4;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_A5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_A6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_AMUX;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_AO5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_AO6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_AX;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_A_CY;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_A_XOR;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_B;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_B1;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_B2;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_B3;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_B4;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_B5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_B6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_BO5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_BO6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_B_CY;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_B_XOR;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_C;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_C1;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_C2;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_C3;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_C4;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_C5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_C6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_CMUX;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_CO5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_CO6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_CX;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_C_CY;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_C_XOR;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_D;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_D1;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_D2;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_D3;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_D4;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_D5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_D6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_DO5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_DO6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_D_CY;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_D_XOR;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X110Y120_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_A;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_A1;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_A2;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_A3;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_A4;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_A5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_A6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_AMUX;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_AO5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_AO6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_AX;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_A_CY;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_A_XOR;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_B;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_B1;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_B2;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_B3;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_B4;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_B5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_B6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_BO5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_BO6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_B_CY;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_B_XOR;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_C;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_C1;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_C2;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_C3;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_C4;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_C5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_C6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_CO5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_CO6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_C_CY;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_C_XOR;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_D;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_D1;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_D2;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_D3;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_D4;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_D5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_D6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_DO5;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_DO6;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_D_CY;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_D_XOR;
  wire [0:0] CLBLL_R_X73Y120_SLICE_X111Y120_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_AMUX;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_AO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_AO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_AX;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_A_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_BO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_BO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_B_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_CO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_CO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_C_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_DO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_DO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_D_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X110Y121_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_AMUX;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_AO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_AO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_AX;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_A_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_BO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_BO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_B_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_CMUX;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_CO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_CO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_CX;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_C_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D1;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D2;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D3;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D4;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_DO5;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_DO6;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D_CY;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_D_XOR;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y121_SLICE_X111Y121_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_AO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_AO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_A_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_BO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_BO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_B_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_CO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_CO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_C_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_DO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_DO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X110Y122_D_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_AO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_AO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_A_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_BO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_BO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_B_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_CO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_CO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_C_XOR;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D1;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D2;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D3;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D4;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_DO5;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_DO6;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D_CY;
  wire [0:0] CLBLL_R_X73Y122_SLICE_X111Y122_D_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_AMUX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_AO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_AO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_AX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_A_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_BO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_BO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_B_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_CO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_CO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_C_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_DO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_DO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_D_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X110Y123_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_AO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_AO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_AX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_A_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_BMUX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_BO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_BO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_BX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_B_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_CO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_CO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_CX;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_C_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D1;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D2;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D3;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D4;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_DO5;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_DO6;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D_CY;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_D_XOR;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y123_SLICE_X111Y123_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_AO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_AO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_AX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_A_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_BMUX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_BO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_BO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_BX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_B_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_CO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_CO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_CX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_C_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_DO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_DO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_D_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X110Y124_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_AMUX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_AO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_AO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_AX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_A_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_BO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_BO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_B_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_CMUX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_CO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_CO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_CX;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_C_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D1;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D2;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D3;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D4;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_DO5;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_DO6;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D_CY;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_D_XOR;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y124_SLICE_X111Y124_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_AO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_AO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_AX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_A_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_BMUX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_BO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_BO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_BX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_B_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_CO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_CO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_CX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_C_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_DO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_DO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_D_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X110Y125_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_AO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_AO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_AX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_A_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_BMUX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_BO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_BO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_BX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_B_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_CO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_CO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_CX;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_C_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D1;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D2;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D3;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D4;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_DO5;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_DO6;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D_CY;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_D_XOR;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y125_SLICE_X111Y125_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_AO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_AO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_AX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_A_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_BMUX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_BO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_BO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_BX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_B_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_CO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_CO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_CX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_C_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_DO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_DO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_D_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X110Y126_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_AMUX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_AO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_AO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_AX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_A_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_BO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_BO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_B_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_CMUX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_CO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_CO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_CX;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_C_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D1;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D2;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D3;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D4;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_DO5;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_DO6;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D_CY;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_D_XOR;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y126_SLICE_X111Y126_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_AO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_AO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_AX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_A_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_BMUX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_BO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_BO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_BX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_B_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_CO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_CO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_CX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_C_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_DO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_DO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_D_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X110Y127_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_AMUX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_AO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_AO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_AX;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_A_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_BO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_BO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_B_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_CO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_CO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_C_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D1;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D2;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D3;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D4;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_DO5;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_DO6;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D_CY;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_D_XOR;
  wire [0:0] CLBLL_R_X73Y127_SLICE_X111Y127_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_AO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_AO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_AX;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_A_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_BMUX;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_BO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_BO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_BX;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_B_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_CO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_CO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_CX;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_C_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_DO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_DO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_D_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X110Y128_F8MUX_O;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_AMUX;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_AO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_AO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_AX;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_A_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_BO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_BO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_B_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_CMUX;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_CO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_CO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_CX;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_C_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D1;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D2;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D3;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D4;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_DO5;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_DO6;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D_CY;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_D_XOR;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y128_SLICE_X111Y128_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_A;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_A1;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_A2;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_A3;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_A4;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_A5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_A6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_AMUX;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_AO5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_AO6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_AX;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_A_CY;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_A_XOR;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_B;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_B1;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_B2;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_B3;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_B4;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_B5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_B6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_BO5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_BO6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_B_CY;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_B_XOR;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_C;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_C1;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_C2;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_C3;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_C4;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_C5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_C6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_CO5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_CO6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_C_CY;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_C_XOR;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_D;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_D1;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_D2;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_D3;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_D4;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_D5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_D6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_DO5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_DO6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_D_CY;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_D_XOR;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X110Y129_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_A;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_A1;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_A2;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_A3;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_A4;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_A5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_A6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_AO5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_AO6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_AX;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_A_CY;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_A_XOR;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_B;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_B1;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_B2;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_B3;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_B4;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_B5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_B6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_BMUX;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_BO5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_BO6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_BX;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_B_CY;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_B_XOR;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_C;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_C1;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_C2;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_C3;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_C4;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_C5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_C6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_CO5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_CO6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_CX;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_C_CY;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_C_XOR;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_D;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_D1;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_D2;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_D3;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_D4;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_D5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_D6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_DO5;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_DO6;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_D_CY;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_D_XOR;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_F7AMUX_O;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_F7BMUX_O;
  wire [0:0] CLBLL_R_X73Y129_SLICE_X111Y129_F8MUX_O;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_A;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_A1;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_A2;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_A3;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_A4;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_A5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_A6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_AMUX;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_AO5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_AO6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_AX;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_A_CY;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_A_XOR;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_B;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_B1;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_B2;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_B3;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_B4;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_B5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_B6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_BO5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_BO6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_B_CY;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_B_XOR;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_C;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_C1;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_C2;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_C3;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_C4;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_C5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_C6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_CO5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_CO6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_C_CY;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_C_XOR;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_D;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_D1;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_D2;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_D3;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_D4;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_D5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_D6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_DO5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_DO6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_D_CY;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_D_XOR;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X114Y115_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_A;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_A1;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_A2;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_A3;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_A4;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_A5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_A6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_AO5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_AO6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_AX;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_A_CY;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_A_XOR;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_B;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_B1;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_B2;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_B3;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_B4;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_B5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_B6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_BMUX;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_BO5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_BO6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_BX;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_B_CY;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_B_XOR;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_C;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_C1;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_C2;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_C3;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_C4;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_C5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_C6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_CO5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_CO6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_CX;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_C_CY;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_C_XOR;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_D;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_D1;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_D2;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_D3;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_D4;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_D5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_D6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_DO5;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_DO6;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_D_CY;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_D_XOR;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y115_SLICE_X115Y115_F8MUX_O;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_A;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_A1;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_A2;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_A3;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_A4;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_A5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_A6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_AMUX;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_AO5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_AO6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_AX;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_A_CY;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_A_XOR;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_B;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_B1;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_B2;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_B3;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_B4;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_B5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_B6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_BO5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_BO6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_B_CY;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_B_XOR;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_C;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_C1;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_C2;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_C3;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_C4;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_C5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_C6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_CO5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_CO6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_C_CY;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_C_XOR;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_D;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_D1;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_D2;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_D3;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_D4;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_D5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_D6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_DO5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_DO6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_D_CY;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_D_XOR;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X114Y116_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_A;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_A1;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_A2;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_A3;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_A4;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_A5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_A6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_AMUX;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_AO5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_AO6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_AX;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_A_CY;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_A_XOR;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_B;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_B1;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_B2;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_B3;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_B4;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_B5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_B6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_BO5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_BO6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_B_CY;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_B_XOR;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_C;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_C1;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_C2;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_C3;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_C4;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_C5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_C6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_CO5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_CO6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_C_CY;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_C_XOR;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_D;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_D1;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_D2;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_D3;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_D4;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_D5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_D6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_DO5;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_DO6;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_D_CY;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_D_XOR;
  wire [0:0] CLBLL_R_X75Y116_SLICE_X115Y116_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_A;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_A1;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_A2;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_A3;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_A4;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_A5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_A6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_AMUX;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_AO5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_AO6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_AX;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_A_CY;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_A_XOR;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_B;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_B1;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_B2;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_B3;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_B4;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_B5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_B6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_BO5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_BO6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_B_CY;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_B_XOR;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_C;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_C1;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_C2;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_C3;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_C4;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_C5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_C6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_CMUX;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_CO5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_CO6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_CX;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_C_CY;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_C_XOR;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_D;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_D1;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_D2;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_D3;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_D4;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_D5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_D6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_DO5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_DO6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_D_CY;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_D_XOR;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X114Y117_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_A;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_A1;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_A2;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_A3;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_A4;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_A5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_A6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_AO5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_AO6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_AX;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_A_CY;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_A_XOR;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_B;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_B1;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_B2;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_B3;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_B4;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_B5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_B6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_BMUX;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_BO5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_BO6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_BX;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_B_CY;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_B_XOR;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_C;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_C1;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_C2;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_C3;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_C4;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_C5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_C6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_CO5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_CO6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_CX;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_C_CY;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_C_XOR;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_D;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_D1;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_D2;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_D3;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_D4;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_D5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_D6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_DO5;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_DO6;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_D_CY;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_D_XOR;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y117_SLICE_X115Y117_F8MUX_O;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_A;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_A1;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_A2;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_A3;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_A4;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_A5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_A6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_AMUX;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_AO5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_AO6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_AX;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_A_CY;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_A_XOR;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_B;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_B1;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_B2;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_B3;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_B4;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_B5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_B6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_BO5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_BO6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_B_CY;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_B_XOR;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_C;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_C1;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_C2;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_C3;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_C4;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_C5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_C6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_CO5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_CO6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_C_CY;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_C_XOR;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_D;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_D1;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_D2;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_D3;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_D4;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_D5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_D6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_DO5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_D_CY;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_D_XOR;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X114Y118_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_A;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_A1;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_A2;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_A3;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_A4;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_A5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_A6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_AO5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_AO6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_AX;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_A_CY;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_A_XOR;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_B;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_B1;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_B2;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_B3;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_B4;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_B5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_B6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_BMUX;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_BO5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_BO6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_BX;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_B_CY;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_B_XOR;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_C;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_C1;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_C2;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_C3;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_C4;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_C5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_C6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_CO5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_CO6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_CX;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_C_CY;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_C_XOR;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_D;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_D1;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_D2;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_D3;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_D4;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_D5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_D6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_DO5;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_DO6;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_D_CY;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_D_XOR;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y118_SLICE_X115Y118_F8MUX_O;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_A;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_A1;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_A2;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_A3;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_A4;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_A5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_A6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_AMUX;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_AO5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_AO6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_AX;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_A_CY;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_A_XOR;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_B;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_B1;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_B2;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_B3;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_B4;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_B5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_B6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_BO5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_BO6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_B_CY;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_B_XOR;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_C;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_C1;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_C2;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_C3;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_C4;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_C5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_C6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_CO5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_CO6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_C_CY;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_C_XOR;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_D;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_D1;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_D2;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_D3;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_D4;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_D5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_D6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_DO5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_DO6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_D_CY;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_D_XOR;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X114Y119_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_A;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_A1;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_A2;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_A3;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_A4;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_A5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_A6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_AMUX;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_AO5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_AO6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_AX;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_A_CY;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_A_XOR;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_B;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_B1;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_B2;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_B3;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_B4;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_B5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_B6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_BO5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_BO6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_B_CY;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_B_XOR;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_C;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_C1;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_C2;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_C3;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_C4;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_C5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_C6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_CO5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_CO6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_C_CY;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_C_XOR;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_D;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_D1;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_D2;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_D3;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_D4;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_D5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_D6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_DO5;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_DO6;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_D_CY;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_D_XOR;
  wire [0:0] CLBLL_R_X75Y119_SLICE_X115Y119_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_A;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_A1;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_A2;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_A3;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_A4;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_A5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_A6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_AO5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_AO6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_AX;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_A_CY;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_A_XOR;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_B;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_B1;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_B2;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_B3;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_B4;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_B5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_B6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_BMUX;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_BO5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_BO6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_BX;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_B_CY;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_B_XOR;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_C;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_C1;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_C2;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_C3;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_C4;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_C5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_C6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_CO5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_CO6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_CX;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_C_CY;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_C_XOR;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_D;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_D1;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_D2;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_D3;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_D4;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_D5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_D6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_DO5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_DO6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_D_CY;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_D_XOR;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X114Y120_F8MUX_O;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_A;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_A1;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_A2;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_A3;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_A4;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_A5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_A6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_AMUX;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_AO5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_AO6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_AX;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_A_CY;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_A_XOR;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_B;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_B1;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_B2;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_B3;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_B4;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_B5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_B6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_BO5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_BO6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_B_CY;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_B_XOR;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_C;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_C1;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_C2;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_C3;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_C4;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_C5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_C6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_CO5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_CO6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_C_CY;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_C_XOR;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_D;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_D1;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_D2;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_D3;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_D4;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_D5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_D6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_DO5;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_DO6;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_D_CY;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_D_XOR;
  wire [0:0] CLBLL_R_X75Y120_SLICE_X115Y120_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_AO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_A_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_BO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_BO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_B_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_CO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_CO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_C_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_DO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_DO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X114Y123_D_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_AO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_AO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_A_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_BO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_BO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_B_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_CO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_CO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_C_XOR;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D1;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D2;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D3;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D4;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_DO5;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D_CY;
  wire [0:0] CLBLL_R_X75Y123_SLICE_X115Y123_D_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_AO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_AO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_AX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_A_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_BMUX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_BO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_BO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_BX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_B_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_CO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_CO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_CX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_C_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_DO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_DO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_D_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X114Y124_F8MUX_O;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_AMUX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_AO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_AO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_AX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_A_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_BO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_BO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_B_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_CMUX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_CO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_CO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_CX;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_C_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D1;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D2;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D3;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D4;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_DO5;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_DO6;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D_CY;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_D_XOR;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y124_SLICE_X115Y124_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_A;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_A1;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_A2;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_A3;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_A4;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_A5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_A6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_AMUX;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_AO5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_AO6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_AX;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_A_CY;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_A_XOR;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_B;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_B1;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_B2;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_B3;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_B4;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_B5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_B6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_BO5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_BO6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_B_CY;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_B_XOR;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_C;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_C1;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_C2;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_C3;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_C4;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_C5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_C6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_CO5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_CO6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_C_CY;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_C_XOR;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_D;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_D1;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_D2;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_D3;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_D4;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_D5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_D6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_DO5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_DO6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_D_CY;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_D_XOR;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X114Y125_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_A;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_A1;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_A2;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_A3;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_A4;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_A5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_A6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_AMUX;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_AO5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_AO6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_AX;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_A_CY;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_A_XOR;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_B;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_B1;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_B2;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_B3;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_B4;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_B5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_B6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_BO5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_BO6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_B_CY;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_B_XOR;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_C;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_C1;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_C2;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_C3;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_C4;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_C5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_C6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_CO5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_CO6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_C_CY;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_C_XOR;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_D;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_D1;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_D2;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_D3;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_D4;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_D5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_D6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_DO5;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_DO6;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_D_CY;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_D_XOR;
  wire [0:0] CLBLL_R_X75Y125_SLICE_X115Y125_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_A;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_A1;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_A2;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_A3;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_A4;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_A5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_A6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_AO5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_AO6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_A_CY;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_A_XOR;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_B;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_B1;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_B2;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_B3;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_B4;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_B5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_B6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_BO5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_BO6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_B_CY;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_B_XOR;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_C;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_C1;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_C2;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_C3;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_C4;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_C5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_C6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_CO5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_CO6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_C_CY;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_C_XOR;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_D;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_D1;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_D2;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_D3;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_D4;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_D5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_D6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_DO5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_DO6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_D_CY;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X114Y126_D_XOR;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_A;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_A1;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_A2;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_A3;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_A4;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_A5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_A6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_AMUX;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_AO5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_AO6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_AX;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_A_CY;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_A_XOR;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_B;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_B1;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_B2;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_B3;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_B4;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_B5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_B6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_BO5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_BO6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_B_CY;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_B_XOR;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_C;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_C1;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_C2;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_C3;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_C4;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_C5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_C6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_CMUX;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_CO5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_CO6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_CX;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_C_CY;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_C_XOR;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_D;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_D1;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_D2;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_D3;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_D4;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_D5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_D6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_DO5;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_DO6;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_D_CY;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_D_XOR;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y126_SLICE_X115Y126_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_AMUX;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_AO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_AO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_AX;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_A_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_BO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_BO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_B_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_CO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_CO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_C_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_DO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_DO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_D_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X114Y127_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_AO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_AO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_AX;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_A_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_BMUX;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_BO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_BO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_BX;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_B_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_CO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_CO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_CX;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_C_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D1;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D2;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D3;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D4;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_DO5;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_DO6;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D_CY;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_D_XOR;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y127_SLICE_X115Y127_F8MUX_O;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_AO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_AX;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_A_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_BMUX;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_BO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_BX;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_B_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_CO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_CO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_CX;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_C_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_DO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_D_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_F7AMUX_O;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_F7BMUX_O;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X114Y128_F8MUX_O;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_AMUX;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_AO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_AX;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_A_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_BO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_B_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_CO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_C_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D1;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D2;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D3;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D4;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_DO5;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D_CY;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_D_XOR;
  wire [0:0] CLBLL_R_X75Y128_SLICE_X115Y128_F7AMUX_O;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_AO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_A_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_BO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_B_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_CO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_C_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_DO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X118Y113_D_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_AO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_AO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_A_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_BO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_BO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_B_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_CO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_CO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_C_XOR;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D1;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D2;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D3;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D4;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_DO5;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_DO6;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D_CY;
  wire [0:0] CLBLL_R_X77Y113_SLICE_X119Y113_D_XOR;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_A;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_A1;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_A2;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_A3;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_A4;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_A5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_A6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_AO5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_A_CY;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_A_XOR;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_B;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_B1;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_B2;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_B3;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_B4;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_B5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_B6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_BO5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_B_CY;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_B_XOR;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_C;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_C1;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_C2;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_C3;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_C4;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_C5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_C6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_CO5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_CO6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_C_CY;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_C_XOR;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_D;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_D1;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_D2;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_D3;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_D4;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_D5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_D6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_DO5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_DO6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_D_CY;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X118Y114_D_XOR;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_A;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_A1;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_A2;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_A3;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_A4;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_A5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_A6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_AO5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_AO6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_A_CY;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_A_XOR;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_B;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_B1;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_B2;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_B3;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_B4;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_B5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_B6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_BO5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_BO6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_B_CY;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_B_XOR;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_C;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_C1;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_C2;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_C3;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_C4;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_C5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_C6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_CO5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_CO6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_C_CY;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_C_XOR;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_D;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_D1;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_D2;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_D3;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_D4;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_D5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_D6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_DO5;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_DO6;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_D_CY;
  wire [0:0] CLBLL_R_X77Y114_SLICE_X119Y114_D_XOR;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_A;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_A1;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_A2;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_A3;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_A4;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_A5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_A6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_AO5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_A_CY;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_A_XOR;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_B;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_B1;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_B2;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_B3;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_B4;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_B5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_B6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_BO5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_BO6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_B_CY;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_B_XOR;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_C;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_C1;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_C2;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_C3;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_C4;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_C5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_C6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_CO5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_CO6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_C_CY;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_C_XOR;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_D;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_D1;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_D2;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_D3;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_D4;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_D5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_D6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_DO5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_DO6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_D_CY;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X118Y115_D_XOR;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_A;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_A1;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_A2;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_A3;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_A4;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_A5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_A6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_AO5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_AO6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_A_CY;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_A_XOR;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_B;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_B1;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_B2;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_B3;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_B4;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_B5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_B6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_BO5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_BO6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_B_CY;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_B_XOR;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_C;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_C1;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_C2;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_C3;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_C4;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_C5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_C6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_CO5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_CO6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_C_CY;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_C_XOR;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_D;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_D1;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_D2;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_D3;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_D4;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_D5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_D6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_DO5;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_DO6;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_D_CY;
  wire [0:0] CLBLL_R_X77Y115_SLICE_X119Y115_D_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_AO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_A_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_BO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_B_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_CO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_C_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_DO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X118Y122_D_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_AO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_AO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_A_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_BO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_BO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_B_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_CO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_CO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_C_XOR;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D1;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D2;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D3;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D4;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_DO5;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_DO6;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D_CY;
  wire [0:0] CLBLL_R_X77Y122_SLICE_X119Y122_D_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_AO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_AO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_AX;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_A_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_BMUX;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_BO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_BO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_BX;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_B_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_CO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_CO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_CX;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_C_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_DO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_DO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_D_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_F7AMUX_O;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_F7BMUX_O;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X118Y125_F8MUX_O;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_AO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_AO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_A_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_BO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_BO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_B_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_CO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_CO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_C_XOR;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D1;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D2;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D3;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D4;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_DO5;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_DO6;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D_CY;
  wire [0:0] CLBLL_R_X77Y125_SLICE_X119Y125_D_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_AO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_A_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_BO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_B_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_CO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_C_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_DO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X118Y129_D_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_AO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_AO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_A_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_BO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_BO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_B_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_CO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_CO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_C_XOR;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D1;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D2;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D3;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D4;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_DO5;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_DO6;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D_CY;
  wire [0:0] CLBLL_R_X77Y129_SLICE_X119Y129_D_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_AO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_A_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_BO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_B_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_CO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_C_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_DO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X118Y130_D_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_AO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_AO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_A_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_BO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_BO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_B_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_CO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_CO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_C_XOR;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D1;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D2;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D3;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D4;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_DO5;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_DO6;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D_CY;
  wire [0:0] CLBLL_R_X77Y130_SLICE_X119Y130_D_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_AO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_A_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_BO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_B_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_CO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_C_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_DO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X118Y131_D_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_AO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_AO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_A_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_BO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_BO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_B_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_CO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_CO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_C_XOR;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D1;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D2;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D3;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D4;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_DO5;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_DO6;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D_CY;
  wire [0:0] CLBLL_R_X77Y131_SLICE_X119Y131_D_XOR;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_A;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_A1;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_A2;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_A3;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_A4;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_A5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_A6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_AO5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_A_CY;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_A_XOR;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_B;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_B1;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_B2;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_B3;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_B4;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_B5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_B6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_BO5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_B_CY;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_B_XOR;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_C;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_C1;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_C2;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_C3;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_C4;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_C5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_C6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_CO5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_CO6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_C_CY;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_C_XOR;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_D;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_D1;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_D2;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_D3;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_D4;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_D5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_D6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_DO5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_DO6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_D_CY;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X118Y133_D_XOR;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_A;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_A1;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_A2;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_A3;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_A4;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_A5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_A6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_AO5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_AO6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_A_CY;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_A_XOR;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_B;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_B1;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_B2;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_B3;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_B4;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_B5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_B6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_BO5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_BO6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_B_CY;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_B_XOR;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_C;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_C1;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_C2;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_C3;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_C4;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_C5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_C6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_CO5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_CO6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_C_CY;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_C_XOR;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_D;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_D1;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_D2;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_D3;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_D4;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_D5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_D6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_DO5;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_DO6;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_D_CY;
  wire [0:0] CLBLL_R_X77Y133_SLICE_X119Y133_D_XOR;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_A;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_A1;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_A2;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_A3;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_A4;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_A5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_A6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_AO5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_A_CY;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_A_XOR;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_B;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_B1;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_B2;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_B3;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_B4;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_B5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_B6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_BO5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_B_CY;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_B_XOR;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_C;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_C1;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_C2;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_C3;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_C4;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_C5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_C6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_CO5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_CO6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_C_CY;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_C_XOR;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_D;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_D1;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_D2;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_D3;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_D4;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_D5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_D6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_DO5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_DO6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_D_CY;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X122Y123_D_XOR;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_A;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_A1;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_A2;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_A3;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_A4;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_A5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_A6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_AO5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_AO6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_A_CY;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_A_XOR;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_B;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_B1;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_B2;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_B3;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_B4;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_B5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_B6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_BO5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_BO6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_B_CY;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_B_XOR;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_C;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_C1;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_C2;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_C3;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_C4;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_C5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_C6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_CO5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_CO6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_C_CY;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_C_XOR;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_D;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_D1;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_D2;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_D3;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_D4;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_D5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_D6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_DO5;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_DO6;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_D_CY;
  wire [0:0] CLBLL_R_X79Y123_SLICE_X123Y123_D_XOR;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_A;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_A1;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_A2;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_A3;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_A4;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_A5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_A6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_AO5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_A_CY;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_A_XOR;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_B;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_B1;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_B2;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_B3;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_B4;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_B5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_B6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_BO5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_B_CY;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_B_XOR;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_C;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_C1;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_C2;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_C3;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_C4;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_C5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_C6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_CO5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_C_CY;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_C_XOR;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_D;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_D1;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_D2;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_D3;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_D4;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_D5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_D6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_DO5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_DO6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_D_CY;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X122Y124_D_XOR;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_A;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_A1;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_A2;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_A3;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_A4;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_A5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_A6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_AO5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_AO6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_A_CY;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_A_XOR;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_B;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_B1;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_B2;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_B3;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_B4;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_B5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_B6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_BO5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_BO6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_B_CY;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_B_XOR;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_C;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_C1;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_C2;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_C3;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_C4;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_C5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_C6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_CO5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_CO6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_C_CY;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_C_XOR;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_D;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_D1;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_D2;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_D3;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_D4;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_D5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_D6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_DO5;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_DO6;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_D_CY;
  wire [0:0] CLBLL_R_X79Y124_SLICE_X123Y124_D_XOR;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_A;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_A1;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_A2;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_A3;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_A4;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_A5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_A6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_AO5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_A_CY;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_A_XOR;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_B;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_B1;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_B2;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_B3;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_B4;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_B5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_B6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_BO5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_BO6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_B_CY;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_B_XOR;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_C;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_C1;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_C2;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_C3;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_C4;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_C5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_C6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_CO5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_CO6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_C_CY;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_C_XOR;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_D;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_D1;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_D2;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_D3;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_D4;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_D5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_D6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_DO5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_DO6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_D_CY;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X122Y125_D_XOR;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_A;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_A1;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_A2;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_A3;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_A4;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_A5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_A6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_AO5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_AO6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_A_CY;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_A_XOR;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_B;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_B1;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_B2;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_B3;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_B4;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_B5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_B6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_BO5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_BO6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_B_CY;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_B_XOR;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_C;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_C1;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_C2;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_C3;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_C4;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_C5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_C6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_CO5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_CO6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_C_CY;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_C_XOR;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_D;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_D1;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_D2;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_D3;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_D4;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_D5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_D6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_DO5;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_DO6;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_D_CY;
  wire [0:0] CLBLL_R_X79Y125_SLICE_X123Y125_D_XOR;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_A;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_A1;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_A2;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_A3;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_A4;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_A5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_A6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_AO5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_A_CY;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_A_XOR;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_B;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_B1;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_B2;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_B3;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_B4;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_B5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_B6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_BO5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_BO6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_B_CY;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_B_XOR;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_C;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_C1;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_C2;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_C3;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_C4;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_C5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_C6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_CO5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_CO6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_C_CY;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_C_XOR;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_D;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_D1;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_D2;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_D3;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_D4;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_D5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_D6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_DO5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_DO6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_D_CY;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X66Y118_D_XOR;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_A;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_A1;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_A2;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_A3;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_A4;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_A5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_A6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_AO5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_AO6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_A_CY;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_A_XOR;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_B;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_B1;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_B2;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_B3;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_B4;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_B5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_B6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_BO5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_BO6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_B_CY;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_B_XOR;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_C;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_C1;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_C2;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_C3;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_C4;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_C5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_C6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_CO5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_CO6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_C_CY;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_C_XOR;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_D;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_D1;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_D2;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_D3;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_D4;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_D5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_D6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_DO5;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_DO6;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_D_CY;
  wire [0:0] CLBLM_L_X44Y118_SLICE_X67Y118_D_XOR;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_A;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_A1;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_A2;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_A3;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_A4;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_A5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_A6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_AO5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_A_CY;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_A_XOR;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_B;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_B1;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_B2;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_B3;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_B4;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_B5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_B6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_BO5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_B_CY;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_B_XOR;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_C;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_C1;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_C2;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_C3;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_C4;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_C5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_C6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_CO5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_CO6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_C_CY;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_C_XOR;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_D;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_D1;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_D2;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_D3;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_D4;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_D5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_D6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_DO5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_DO6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_D_CY;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X70Y116_D_XOR;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_A;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_A1;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_A2;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_A3;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_A4;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_A5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_A6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_AO5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_AO6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_A_CY;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_A_XOR;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_B;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_B1;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_B2;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_B3;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_B4;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_B5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_B6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_BO5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_BO6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_B_CY;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_B_XOR;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_C;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_C1;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_C2;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_C3;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_C4;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_C5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_C6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_CO5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_CO6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_C_CY;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_C_XOR;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_D;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_D1;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_D2;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_D3;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_D4;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_D5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_D6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_DO5;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_DO6;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_D_CY;
  wire [0:0] CLBLM_L_X46Y116_SLICE_X71Y116_D_XOR;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_A;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_A1;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_A2;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_A3;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_A4;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_A5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_A6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_AMUX;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_AO5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_AO6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_AQ;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_AX;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_A_CY;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_A_XOR;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_B;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_B1;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_B2;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_B3;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_B4;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_B5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_B6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_BO5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_BO6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_BQ;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_BX;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_B_CY;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_B_XOR;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_C;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_C1;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_C2;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_C3;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_C4;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_C5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_C6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_CLK;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_CMUX;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_CO5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_CO6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_C_CY;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_C_XOR;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_D;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_D1;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_D2;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_D3;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_D4;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_D5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_D6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_DO5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_DO6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_D_CY;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X84Y116_D_XOR;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_A;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_A1;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_A2;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_A3;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_A4;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_A5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_A6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_AO5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_AO6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_A_CY;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_A_XOR;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_B;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_B1;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_B2;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_B3;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_B4;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_B5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_B6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_BO5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_BO6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_B_CY;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_B_XOR;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_C;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_C1;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_C2;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_C3;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_C4;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_C5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_C6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_CO5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_CO6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_C_CY;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_C_XOR;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_D;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_D1;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_D2;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_D3;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_D4;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_D5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_D6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_DO5;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_DO6;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_D_CY;
  wire [0:0] CLBLM_L_X56Y116_SLICE_X85Y116_D_XOR;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_A;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_A1;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_A2;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_A3;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_A4;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_A5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_A6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_AO5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_AO6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_A_CY;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_A_XOR;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_B;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_B1;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_B2;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_B3;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_B4;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_B5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_B6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_BO5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_BO6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_B_CY;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_B_XOR;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_C;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_C1;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_C2;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_C3;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_C4;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_C5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_C6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_CO5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_CO6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_C_CY;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_C_XOR;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_D;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_D1;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_D2;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_D3;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_D4;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_D5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_D6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_DO5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_DO6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_D_CY;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X102Y119_D_XOR;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_A;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_A1;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_A2;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_A3;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_A4;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_A5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_A6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_AO5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_AO6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_A_CY;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_A_XOR;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_B;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_B1;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_B2;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_B3;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_B4;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_B5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_B6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_BO5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_BO6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_B_CY;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_B_XOR;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_C;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_C1;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_C2;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_C3;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_C4;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_C5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_C6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_CO5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_CO6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_C_CY;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_C_XOR;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_D;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_D1;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_D2;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_D3;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_D4;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_D5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_D6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_DO5;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_DO6;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_D_CY;
  wire [0:0] CLBLM_L_X68Y119_SLICE_X103Y119_D_XOR;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_A;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_A1;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_A2;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_A3;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_A4;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_A5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_A6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_AO5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_AO6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_A_CY;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_A_XOR;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_B;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_B1;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_B2;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_B3;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_B4;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_B5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_B6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_BO5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_BO6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_B_CY;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_B_XOR;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_C;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_C1;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_C2;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_C3;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_C4;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_C5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_C6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_CO5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_CO6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_C_CY;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_C_XOR;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_D;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_D1;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_D2;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_D3;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_D4;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_D5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_D6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_DO5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_DO6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_D_CY;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X104Y117_D_XOR;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_A;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_A1;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_A2;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_A3;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_A4;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_A5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_A6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_AO5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_AO6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_A_CY;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_A_XOR;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_B;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_B1;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_B2;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_B3;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_B4;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_B5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_B6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_BO5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_BO6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_B_CY;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_B_XOR;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_C;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_C1;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_C2;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_C3;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_C4;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_C5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_C6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_CO5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_CO6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_C_CY;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_C_XOR;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_D;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_D1;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_D2;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_D3;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_D4;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_D5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_D6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_DO5;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_DO6;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_D_CY;
  wire [0:0] CLBLM_L_X70Y117_SLICE_X105Y117_D_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_AO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_AO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_AQ;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_A_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_BMUX;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_BO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_BO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_B_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_CLK;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_CO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_CO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_C_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_DO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_DO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X104Y119_D_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_AO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_AO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_AX;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_A_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_BO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_BO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_BQ;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_BX;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_B_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_CLK;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_CO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_C_XOR;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D1;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D2;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D3;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D4;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_DO5;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_DO6;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D_CY;
  wire [0:0] CLBLM_L_X70Y119_SLICE_X105Y119_D_XOR;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_A;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_A1;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_A2;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_A3;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_A4;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_A5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_A6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_AO5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_AO6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_AQ;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_AX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_A_CY;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_A_XOR;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_B;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_B1;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_B2;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_B3;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_B4;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_B5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_B6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_BMUX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_BO5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_BO6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_BQ;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_BX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_B_CY;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_B_XOR;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_C;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_C1;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_C2;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_C3;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_C4;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_C5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_C6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_CLK;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_CMUX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_CO5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_CO6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_CQ;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_CX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_C_CY;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_C_XOR;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_D;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_D1;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_D2;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_D3;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_D4;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_D5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_D6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_DO5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_DO6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_DQ;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_DX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_D_CY;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X104Y121_D_XOR;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_A;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_A1;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_A2;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_A3;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_A4;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_A5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_A6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_AMUX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_AO5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_AO6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_AQ;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_AX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_A_CY;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_A_XOR;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_B;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_B1;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_B2;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_B3;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_B4;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_B5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_B6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_BMUX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_BO5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_BO6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_BQ;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_BX;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_B_CY;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_B_XOR;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_C;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_C1;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_C2;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_C3;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_C4;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_C5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_C6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_CLK;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_CO5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_CO6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_C_CY;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_C_XOR;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_D;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_D1;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_D2;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_D3;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_D4;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_D5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_D6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_DO5;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_DO6;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_D_CY;
  wire [0:0] CLBLM_L_X70Y121_SLICE_X105Y121_D_XOR;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_A;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_A1;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_A2;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_A3;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_A4;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_A5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_A6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_AMUX;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_AO5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_AO6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_AQ;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_AX;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_A_CY;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_A_XOR;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_B;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_B1;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_B2;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_B3;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_B4;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_B5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_B6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_BO5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_BO6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_BQ;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_BX;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_B_CY;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_B_XOR;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_C;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_C1;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_C2;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_C3;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_C4;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_C5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_C6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_CLK;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_CMUX;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_CO5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_CO6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_C_CY;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_C_XOR;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_D;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_D1;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_D2;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_D3;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_D4;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_D5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_D6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_DO5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_DO6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_D_CY;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X104Y122_D_XOR;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_A;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_A1;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_A2;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_A3;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_A4;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_A5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_A6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_AO5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_AO6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_A_CY;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_A_XOR;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_B;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_B1;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_B2;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_B3;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_B4;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_B5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_B6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_BO5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_BO6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_B_CY;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_B_XOR;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_C;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_C1;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_C2;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_C3;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_C4;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_C5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_C6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_CO5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_CO6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_C_CY;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_C_XOR;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_D;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_D1;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_D2;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_D3;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_D4;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_D5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_D6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_DO5;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_DO6;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_D_CY;
  wire [0:0] CLBLM_L_X70Y122_SLICE_X105Y122_D_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_AO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_AO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_A_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_BO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_BO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_B_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_CO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_CO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_C_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_DO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_DO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X104Y123_D_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_AO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_AO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_AQ;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_AX;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_A_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_BO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_BO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_BQ;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_BX;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_B_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_CLK;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_CO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_CQ;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_CX;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_C_XOR;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D1;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D2;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D3;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D4;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_DO5;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_DO6;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D_CY;
  wire [0:0] CLBLM_L_X70Y123_SLICE_X105Y123_D_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_AO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_AO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_AQ;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_AX;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_A_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_BO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_BO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_BQ;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_BX;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_B_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_CLK;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_CO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_CO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_C_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_DO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_DO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X104Y124_D_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_AO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_AQ;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_AX;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_A_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_BO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_B_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_CLK;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_CO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_CO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_C_XOR;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D1;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D2;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D3;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D4;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_DO5;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_DO6;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D_CY;
  wire [0:0] CLBLM_L_X70Y124_SLICE_X105Y124_D_XOR;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_A;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_A1;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_A2;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_A3;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_A4;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_A5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_A6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_AMUX;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_AO5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_AO6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_AQ;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_AX;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_A_CY;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_A_XOR;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_B;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_B1;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_B2;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_B3;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_B4;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_B5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_B6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_BMUX;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_BO5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_BO6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_BQ;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_BX;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_B_CY;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_B_XOR;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_C;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_C1;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_C2;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_C3;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_C4;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_C5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_C6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_CLK;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_CO5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_CO6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_CQ;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_CX;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_C_CY;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_C_XOR;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_D;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_D1;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_D2;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_D3;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_D4;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_D5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_D6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_DO5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_DO6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_D_CY;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X104Y127_D_XOR;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_A;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_A1;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_A2;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_A3;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_A4;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_A5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_A6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_AO5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_AO6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_A_CY;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_A_XOR;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_B;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_B1;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_B2;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_B3;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_B4;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_B5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_B6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_BO5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_BO6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_B_CY;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_B_XOR;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_C;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_C1;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_C2;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_C3;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_C4;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_C5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_C6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_CO5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_CO6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_C_CY;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_C_XOR;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_D;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_D1;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_D2;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_D3;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_D4;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_D5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_D6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_DO5;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_DO6;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_D_CY;
  wire [0:0] CLBLM_L_X70Y127_SLICE_X105Y127_D_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_AO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_AO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_AX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_A_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_BMUX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_BO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_B_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_CLK;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_CO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_CO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_C_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_DO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_DO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X104Y128_D_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_AMUX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_AO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_AQ;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_AX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_A_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_BO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_BO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_BQ;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_BX;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_B_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_CLK;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_CO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_C_XOR;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D1;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D2;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D3;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D4;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_DO5;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_DO6;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D_CY;
  wire [0:0] CLBLM_L_X70Y128_SLICE_X105Y128_D_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_AMUX;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_AO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_AO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_AX;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_A_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_BMUX;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_BO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_BO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_BQ;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_BX;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_B_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_CLK;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_CMUX;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_CO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_C_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_DO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_DO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X104Y129_D_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_AO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_AO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_A_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_BO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_BO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_B_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_CO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_CO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_C_XOR;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D1;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D2;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D3;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D4;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_DO5;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_DO6;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D_CY;
  wire [0:0] CLBLM_L_X70Y129_SLICE_X105Y129_D_XOR;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_A;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_A1;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_A2;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_A3;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_A4;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_A5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_A6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_AO5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_AO6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_A_CY;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_A_XOR;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_B;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_B1;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_B2;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_B3;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_B4;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_B5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_B6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_BO5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_BO6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_B_CY;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_B_XOR;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_C;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_C1;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_C2;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_C3;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_C4;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_C5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_C6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_CO5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_CO6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_C_CY;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_C_XOR;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_D;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_D1;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_D2;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_D3;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_D4;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_D5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_D6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_DO5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_DO6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_D_CY;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X108Y114_D_XOR;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_A;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_A1;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_A2;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_A3;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_A4;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_A5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_A6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_AMUX;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_AO5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_AO6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_AX;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_A_CY;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_A_XOR;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_B;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_B1;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_B2;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_B3;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_B4;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_B5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_B6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_BO5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_BO6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_B_CY;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_B_XOR;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_C;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_C1;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_C2;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_C3;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_C4;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_C5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_C6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_CO5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_CO6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_C_CY;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_C_XOR;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_D;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_D1;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_D2;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_D3;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_D4;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_D5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_D6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_DO5;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_DO6;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_D_CY;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_D_XOR;
  wire [0:0] CLBLM_L_X72Y114_SLICE_X109Y114_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_A;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_A1;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_A2;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_A3;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_A4;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_A5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_A6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_AO5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_AO6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_AX;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_A_CY;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_A_XOR;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_B;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_B1;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_B2;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_B3;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_B4;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_B5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_B6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_BMUX;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_BO5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_BO6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_BX;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_B_CY;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_B_XOR;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_C;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_C1;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_C2;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_C3;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_C4;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_C5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_C6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_CO5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_CO6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_CX;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_C_CY;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_C_XOR;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_D;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_D1;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_D2;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_D3;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_D4;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_D5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_D6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_DO5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_DO6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_D_CY;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_D_XOR;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X108Y115_F8MUX_O;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_A;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_A1;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_A2;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_A3;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_A4;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_A5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_A6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_AMUX;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_AO5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_AO6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_AX;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_A_CY;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_A_XOR;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_B;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_B1;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_B2;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_B3;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_B4;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_B5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_B6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_BO5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_BO6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_B_CY;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_B_XOR;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_C;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_C1;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_C2;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_C3;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_C4;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_C5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_C6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_CMUX;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_CO5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_CO6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_CX;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_C_CY;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_C_XOR;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_D;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_D1;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_D2;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_D3;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_D4;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_D5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_D6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_DO5;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_DO6;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_D_CY;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_D_XOR;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y115_SLICE_X109Y115_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_AMUX;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_AO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_AO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_AX;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_A_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_BO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_BO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_B_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_CO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_CO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_C_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_DO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_DO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_D_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X108Y116_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_AMUX;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_AO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_AO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_AX;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_A_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_BO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_BO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_B_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_CMUX;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_CO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_CO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_CX;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_C_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D1;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D2;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D3;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D4;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_DO5;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_DO6;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D_CY;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_D_XOR;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y116_SLICE_X109Y116_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_AMUX;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_AO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_AO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_AX;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_A_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_BO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_BO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_B_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_CMUX;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_CO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_CO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_CX;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_C_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_DO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_DO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_D_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X108Y117_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_AMUX;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_AO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_AO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_AX;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_A_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_BO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_BO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_B_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_CO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_CO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_C_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D1;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D2;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D3;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D4;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_DO5;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_DO6;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D_CY;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_D_XOR;
  wire [0:0] CLBLM_L_X72Y117_SLICE_X109Y117_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_AMUX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_AO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_AO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_AX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_A_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_BO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_BO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_B_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_CO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_CO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_C_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_DO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_DO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_D_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X108Y118_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_AMUX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_AO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_AO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_AX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_A_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_BO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_BO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_B_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_CMUX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_CO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_CO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_CX;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_C_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D1;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D2;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D3;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D4;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_DO5;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_DO6;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D_CY;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_D_XOR;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y118_SLICE_X109Y118_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_AMUX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_AO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_AO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_AX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_A_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_BO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_BO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_B_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_CO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_CO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_C_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_DO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_D_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X108Y119_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_AMUX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_AO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_AO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_AX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_A_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_BO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_BO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_B_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_CMUX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_CO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_CO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_CX;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_C_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D1;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D2;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D3;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D4;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_DO5;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_DO6;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D_CY;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_D_XOR;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y119_SLICE_X109Y119_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_AMUX;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_AO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_AO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_AX;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_A_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_BO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_BO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_B_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_CO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_CO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_C_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_DO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_DO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_D_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X108Y120_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_AO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_AO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_AX;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_A_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_BMUX;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_BO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_BO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_BX;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_B_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_CO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_CO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_CX;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_C_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D1;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D2;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D3;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D4;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_DO5;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_DO6;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D_CY;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_D_XOR;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y120_SLICE_X109Y120_F8MUX_O;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_AO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_AO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_AX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_A_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_BMUX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_BO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_BO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_BX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_B_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_CO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_CO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_CX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_C_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_DO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_DO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_D_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X108Y121_F8MUX_O;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_AO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_AO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_AX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_A_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_BMUX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_BO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_BO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_BX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_B_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_CO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_CO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_CX;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_C_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D1;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D2;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D3;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D4;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_DO5;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_DO6;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D_CY;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_D_XOR;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y121_SLICE_X109Y121_F8MUX_O;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_AO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_A_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_BO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_BO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_B_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_CO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_CO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_C_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_DO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_DO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X108Y122_D_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_AO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_AO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_A_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_BO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_BO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_B_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_CO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_CO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_C_XOR;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D1;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D2;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D3;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D4;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_DO5;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_DO6;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D_CY;
  wire [0:0] CLBLM_L_X72Y122_SLICE_X109Y122_D_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_AMUX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_AO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_AO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_AX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_A_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_BO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_BO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_B_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_CMUX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_CO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_CO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_CX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_C_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_DO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_DO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_D_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X108Y123_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_AO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_AO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_AX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_A_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_BMUX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_BO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_BO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_BX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_B_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_CO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_CO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_CX;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_C_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D1;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D2;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D3;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D4;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_DO5;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_DO6;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D_CY;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_D_XOR;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y123_SLICE_X109Y123_F8MUX_O;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_AMUX;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_AO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_AO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_AX;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_A_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_BO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_B_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_CO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_CO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_C_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_DO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_DO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_D_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X108Y124_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_AMUX;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_AO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_AO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_AX;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_A_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_BO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_BO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_B_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_CMUX;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_CO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_CO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_CX;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_C_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D1;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D2;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D3;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D4;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_DO5;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_DO6;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D_CY;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_D_XOR;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y124_SLICE_X109Y124_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_AMUX;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_AO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_AO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_AX;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_A_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_BO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_BO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_B_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_CMUX;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_CO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_CO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_CX;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_C_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_DO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_DO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_D_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X108Y125_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_AO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_AO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_AX;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_A_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_BMUX;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_BO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_BO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_BX;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_B_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_CO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_CO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_CX;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_C_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D1;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D2;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D3;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D4;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_DO5;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_DO6;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D_CY;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_D_XOR;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y125_SLICE_X109Y125_F8MUX_O;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_AO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_AO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_AX;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_A_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_BMUX;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_BO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_BO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_BX;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_B_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_CO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_CX;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_C_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_DO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_DO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_D_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X108Y126_F8MUX_O;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_AMUX;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_AO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_AO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_AX;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_A_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_BO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_BO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_B_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_CMUX;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_CO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_CO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_CX;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_C_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D1;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D2;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D3;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D4;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_DO5;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_DO6;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D_CY;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_D_XOR;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y126_SLICE_X109Y126_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_AMUX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_AO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_AO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_AX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_A_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_BO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_BO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_B_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_CMUX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_CO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_CO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_CX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_C_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_DO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_DO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_D_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X108Y127_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_AO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_AO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_AX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_A_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_BMUX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_BO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_BO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_BX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_B_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_CO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_CO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_CX;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_C_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D1;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D2;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D3;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D4;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_DO5;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_DO6;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D_CY;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_D_XOR;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y127_SLICE_X109Y127_F8MUX_O;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_AMUX;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_AO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_AO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_AX;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_A_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_BO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_BO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_B_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_CO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_CO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_C_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_DO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_DO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_D_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X108Y128_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_AMUX;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_AO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_AO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_AX;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_A_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_BO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_BO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_B_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_CO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_CO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_C_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D1;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D2;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D3;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D4;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_DO5;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_DO6;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D_CY;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_D_XOR;
  wire [0:0] CLBLM_L_X72Y128_SLICE_X109Y128_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_AO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_AO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_AX;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_A_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_BMUX;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_BO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_BO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_BX;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_B_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_CO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_CO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_CX;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_C_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_DO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_DO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_D_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X108Y129_F8MUX_O;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_AMUX;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_AO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_AO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_AX;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_A_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_BO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_BO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_B_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_CMUX;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_CO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_CO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_CX;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_C_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D1;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D2;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D3;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D4;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_DO5;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_DO6;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D_CY;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_D_XOR;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_F7AMUX_O;
  wire [0:0] CLBLM_L_X72Y129_SLICE_X109Y129_F7BMUX_O;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_AO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_AO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_AX;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_A_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_BO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_BO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_B_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_CLK;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_CO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_CO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_C_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_DO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_DO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X108Y131_D_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_AO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_AO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_A_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_BO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_BO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_B_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_CO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_CO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_C_XOR;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D1;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D2;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D3;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D4;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_DO5;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_DO6;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D_CY;
  wire [0:0] CLBLM_L_X72Y131_SLICE_X109Y131_D_XOR;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_A;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_A1;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_A2;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_A3;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_A4;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_A5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_A6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_AO5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_AO6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_A_CY;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_A_XOR;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_B;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_B1;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_B2;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_B3;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_B4;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_B5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_B6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_BO5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_BO6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_B_CY;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_B_XOR;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_C;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_C1;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_C2;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_C3;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_C4;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_C5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_C6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_CO5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_CO6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_C_CY;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_C_XOR;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_D;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_D1;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_D2;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_D3;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_D4;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_D5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_D6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_DO5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_DO6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_D_CY;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X112Y115_D_XOR;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_A;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_A1;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_A2;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_A3;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_A4;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_A5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_A6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_AO5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_AO6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_AX;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_A_CY;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_A_XOR;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_B;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_B1;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_B2;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_B3;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_B4;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_B5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_B6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_BMUX;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_BO5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_BO6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_BX;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_B_CY;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_B_XOR;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_C;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_C1;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_C2;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_C3;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_C4;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_C5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_C6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_CO5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_CO6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_CX;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_C_CY;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_C_XOR;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_D;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_D1;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_D2;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_D3;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_D4;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_D5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_D6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_DO5;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_DO6;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_D_CY;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_D_XOR;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y115_SLICE_X113Y115_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_A;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_A1;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_A2;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_A3;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_A4;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_A5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_A6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_AO5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_AO6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_AX;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_A_CY;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_A_XOR;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_B;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_B1;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_B2;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_B3;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_B4;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_B5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_B6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_BMUX;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_BO5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_BO6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_BX;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_B_CY;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_B_XOR;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_C;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_C1;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_C2;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_C3;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_C4;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_C5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_C6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_CO5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_CO6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_CX;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_C_CY;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_C_XOR;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_D;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_D1;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_D2;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_D3;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_D4;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_D5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_D6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_DO5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_DO6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_D_CY;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_D_XOR;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X112Y116_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_A;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_A1;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_A2;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_A3;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_A4;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_A5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_A6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_AMUX;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_AO5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_AO6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_AX;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_A_CY;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_A_XOR;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_B;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_B1;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_B2;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_B3;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_B4;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_B5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_B6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_BO5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_BO6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_B_CY;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_B_XOR;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_C;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_C1;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_C2;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_C3;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_C4;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_C5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_C6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_CO5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_CO6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_C_CY;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_C_XOR;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_D;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_D1;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_D2;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_D3;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_D4;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_D5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_D6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_DO5;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_DO6;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_D_CY;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_D_XOR;
  wire [0:0] CLBLM_L_X74Y116_SLICE_X113Y116_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_AO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_AO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_AX;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_A_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_BMUX;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_BO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_BO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_BX;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_B_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_CO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_CO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_CX;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_C_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_DO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_DO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_D_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X112Y117_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_AMUX;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_AO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_AO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_AX;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_A_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_BO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_BO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_B_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_CO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_CO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_C_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D1;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D2;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D3;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D4;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_DO5;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_DO6;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D_CY;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_D_XOR;
  wire [0:0] CLBLM_L_X74Y117_SLICE_X113Y117_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_AO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_AO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_A_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_BO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_BO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_B_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_CO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_CO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_C_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_DO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_DO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X112Y118_D_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_AMUX;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_AO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_AO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_AX;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_A_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_BO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_BO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_B_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_CO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_CO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_C_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D1;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D2;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D3;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D4;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_DO5;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_DO6;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D_CY;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_D_XOR;
  wire [0:0] CLBLM_L_X74Y118_SLICE_X113Y118_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_AO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_AO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_AX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_A_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_BMUX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_BO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_BO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_BX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_B_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_CO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_CO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_CX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_C_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_DO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_DO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_D_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X112Y119_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_AMUX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_AO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_AO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_AX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_A_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_BO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_BO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_B_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_CMUX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_CO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_CO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_CX;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_C_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D1;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D2;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D3;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D4;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_DO5;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_DO6;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D_CY;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_D_XOR;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y119_SLICE_X113Y119_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_AO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_AX;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_A_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_BMUX;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_BO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_BO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_BX;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_B_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_CO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_CO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_CX;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_C_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_DO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_DO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_D_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X112Y120_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_AMUX;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_AO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_AO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_A_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_BO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_BO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_B_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_CO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_CO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_C_XOR;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D1;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D2;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D3;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D4;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_DO5;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_DO6;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D_CY;
  wire [0:0] CLBLM_L_X74Y120_SLICE_X113Y120_D_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_AO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_AO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_AX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_A_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_BMUX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_BO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_BO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_BX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_B_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_CO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_CO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_CX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_C_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_DO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_DO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_D_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X112Y121_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_AO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_AO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_AX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_A_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_BMUX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_BO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_BO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_BX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_B_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_CO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_CO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_CX;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_C_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D1;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D2;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D3;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D4;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_DO5;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_DO6;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D_CY;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_D_XOR;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y121_SLICE_X113Y121_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_AMUX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_AO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_AO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_AX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_A_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_BO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_BO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_B_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_CO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_CO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_C_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_DO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_DO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_D_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X112Y123_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_AO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_AO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_AX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_A_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_BMUX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_BO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_BO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_BX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_B_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_CO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_CO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_CX;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_C_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D1;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D2;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D3;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D4;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_DO5;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_DO6;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D_CY;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_D_XOR;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y123_SLICE_X113Y123_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_A;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_A1;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_A2;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_A3;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_A4;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_A5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_A6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_AO5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_AO6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_AX;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_A_CY;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_A_XOR;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_B;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_B1;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_B2;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_B3;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_B4;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_B5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_B6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_BMUX;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_BO5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_BO6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_BX;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_B_CY;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_B_XOR;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_C;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_C1;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_C2;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_C3;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_C4;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_C5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_C6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_CO5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_CO6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_CX;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_C_CY;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_C_XOR;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_D;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_D1;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_D2;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_D3;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_D4;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_D5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_D6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_DO5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_DO6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_D_CY;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_D_XOR;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X112Y124_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_A;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_A1;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_A2;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_A3;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_A4;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_A5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_A6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_AMUX;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_AO5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_AO6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_AX;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_A_CY;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_A_XOR;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_B;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_B1;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_B2;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_B3;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_B4;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_B5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_B6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_BO5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_BO6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_B_CY;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_B_XOR;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_C;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_C1;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_C2;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_C3;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_C4;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_C5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_C6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_CMUX;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_CO5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_CO6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_CX;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_C_CY;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_C_XOR;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_D;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_D1;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_D2;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_D3;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_D4;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_D5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_D6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_DO5;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_DO6;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_D_CY;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_D_XOR;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y124_SLICE_X113Y124_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_AMUX;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_AO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_AO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_AX;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_A_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_BO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_BO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_B_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_CO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_CO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_C_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_DO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_DO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_D_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X112Y125_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_AMUX;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_AO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_AO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_AX;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_A_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_BO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_BO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_B_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_CMUX;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_CO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_CO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_CX;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_C_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D1;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D2;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D3;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D4;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_DO5;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_DO6;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D_CY;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_D_XOR;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y125_SLICE_X113Y125_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_AO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_AO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_AX;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_A_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_BMUX;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_BO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_BO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_BX;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_B_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_CO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_CO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_CX;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_C_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_DO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_DO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_D_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X112Y126_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_AO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_AO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_A_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_BO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_BO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_B_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_CO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_CO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_C_XOR;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D1;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D2;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D3;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D4;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_DO5;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_DO6;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D_CY;
  wire [0:0] CLBLM_L_X74Y126_SLICE_X113Y126_D_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_AMUX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_AO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_AO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_AX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_A_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_BO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_BO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_B_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_CMUX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_CO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_CO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_CX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_C_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_DO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_DO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_D_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X112Y127_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_AMUX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_AO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_AO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_AX;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_A_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_BO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_BO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_B_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_CO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_CO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_C_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D1;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D2;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D3;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D4;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_DO5;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_DO6;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D_CY;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_D_XOR;
  wire [0:0] CLBLM_L_X74Y127_SLICE_X113Y127_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_AMUX;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_AO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_AO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_AX;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_A_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_BO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_BO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_B_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_CO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_CO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_C_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_DO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_DO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_D_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X112Y128_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_AO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_AO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_AX;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_A_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_BMUX;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_BO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_BO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_BX;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_B_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_CO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_CO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_CX;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_C_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D1;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D2;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D3;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D4;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_DO5;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_DO6;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D_CY;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_D_XOR;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_F7BMUX_O;
  wire [0:0] CLBLM_L_X74Y128_SLICE_X113Y128_F8MUX_O;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_AMUX;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_AO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_AO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_AX;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_A_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_BO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_BO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_B_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_CO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_CO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_C_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_DO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_DO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_D_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X112Y129_F7AMUX_O;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_AO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_AO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_A_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_BO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_BO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_B_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_CO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_CO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_C_XOR;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D1;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D2;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D3;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D4;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_DO5;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_DO6;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D_CY;
  wire [0:0] CLBLM_L_X74Y129_SLICE_X113Y129_D_XOR;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_A;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_A1;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_A2;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_A3;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_A4;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_A5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_A6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_AO5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_AO6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_AX;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_A_CY;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_A_XOR;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_B;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_B1;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_B2;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_B3;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_B4;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_B5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_B6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_BMUX;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_BO5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_BO6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_BX;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_B_CY;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_B_XOR;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_C;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_C1;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_C2;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_C3;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_C4;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_C5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_C6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_CO5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_CO6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_CX;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_C_CY;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_C_XOR;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_D;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_D1;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_D2;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_D3;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_D4;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_D5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_D6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_DO5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_DO6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_D_CY;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_D_XOR;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_F7AMUX_O;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_F7BMUX_O;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X116Y120_F8MUX_O;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_A;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_A1;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_A2;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_A3;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_A4;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_A5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_A6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_AO5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_AO6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_A_CY;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_A_XOR;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_B;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_B1;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_B2;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_B3;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_B4;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_B5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_B6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_BO5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_BO6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_B_CY;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_B_XOR;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_C;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_C1;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_C2;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_C3;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_C4;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_C5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_C6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_CO5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_CO6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_C_CY;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_C_XOR;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_D;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_D1;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_D2;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_D3;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_D4;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_D5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_D6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_DO5;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_DO6;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_D_CY;
  wire [0:0] CLBLM_L_X76Y120_SLICE_X117Y120_D_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_AMUX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_AO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_AO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_AX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_A_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_BO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_BO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_B_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CMUX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_CX;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_C_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_DO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_DO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_D_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_F7AMUX_O;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X116Y124_F7BMUX_O;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_AO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_AO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_A_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_BO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_BO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_B_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_CO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_CO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_C_XOR;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D1;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D2;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D3;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D4;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_DO5;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_DO6;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D_CY;
  wire [0:0] CLBLM_L_X76Y124_SLICE_X117Y124_D_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_AO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_AO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_AX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_A_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_BMUX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_BO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_BO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_BX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_B_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_CO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_CO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_CX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_C_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_DO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_DO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_D_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_F7AMUX_O;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_F7BMUX_O;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X116Y125_F8MUX_O;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_AO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_AO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_AX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_A_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_BMUX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_BO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_BO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_BX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_B_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_CO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_CO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_CX;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_C_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D1;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D2;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D3;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D4;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_DO5;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_DO6;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D_CY;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_D_XOR;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_F7AMUX_O;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_F7BMUX_O;
  wire [0:0] CLBLM_L_X76Y125_SLICE_X117Y125_F8MUX_O;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_AMUX;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_AO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_AO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_AX;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_A_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_BO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_BO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_B_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_CO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_C_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_DO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_DO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_D_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X116Y127_F7AMUX_O;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_AO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_AO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_A_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_BO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_BO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_B_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_CO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_CO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_C_XOR;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D1;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D2;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D3;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D4;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_DO5;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_DO6;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D_CY;
  wire [0:0] CLBLM_L_X76Y127_SLICE_X117Y127_D_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_AO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_AO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_AX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_A_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_BMUX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_BO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_BO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_BX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_B_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_CO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_CO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_CX;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_C_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_DO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_DO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_D_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_F7AMUX_O;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_F7BMUX_O;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X116Y128_F8MUX_O;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_AO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_AO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_A_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_BO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_BO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_B_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_CO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_CO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_C_XOR;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D1;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D2;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D3;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D4;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_DO5;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_DO6;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D_CY;
  wire [0:0] CLBLM_L_X76Y128_SLICE_X117Y128_D_XOR;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_A;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_A1;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_A2;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_A3;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_A4;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_A5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_A6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_AO5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_A_CY;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_A_XOR;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_B;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_B1;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_B2;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_B3;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_B4;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_B5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_B6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_BO5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_B_CY;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_B_XOR;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_C;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_C1;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_C2;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_C3;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_C4;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_C5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_C6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_CO5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_CO6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_C_CY;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_C_XOR;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_D;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_D1;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_D2;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_D3;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_D4;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_D5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_D6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_DO5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_DO6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_D_CY;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X116Y131_D_XOR;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_A;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_A1;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_A2;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_A3;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_A4;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_A5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_A6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_AO5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_AO6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_A_CY;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_A_XOR;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_B;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_B1;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_B2;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_B3;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_B4;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_B5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_B6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_BO5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_BO6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_B_CY;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_B_XOR;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_C;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_C1;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_C2;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_C3;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_C4;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_C5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_C6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_CO5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_CO6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_C_CY;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_C_XOR;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_D;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_D1;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_D2;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_D3;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_D4;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_D5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_D6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_DO5;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_DO6;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_D_CY;
  wire [0:0] CLBLM_L_X76Y131_SLICE_X117Y131_D_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_AO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_AO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_A_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_BO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_BO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_B_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_CO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_CO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_C_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_DO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_DO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X116Y133_D_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_AO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_A_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_BO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_BO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_B_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_CO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_CO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_C_XOR;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D1;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D2;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D3;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D4;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_DO5;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_DO6;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D_CY;
  wire [0:0] CLBLM_L_X76Y133_SLICE_X117Y133_D_XOR;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_A;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_A1;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_A2;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_A3;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_A4;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_A5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_A6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_AO5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_A_CY;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_A_XOR;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_B;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_B1;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_B2;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_B3;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_B4;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_B5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_B6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_BO5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_B_CY;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_B_XOR;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_C;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_C1;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_C2;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_C3;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_C4;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_C5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_C6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_CO5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_CO6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_C_CY;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_C_XOR;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_D;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_D1;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_D2;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_D3;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_D4;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_D5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_D6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_DO5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_DO6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_D_CY;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X120Y117_D_XOR;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_A;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_A1;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_A2;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_A3;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_A4;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_A5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_A6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_AO5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_AO6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_A_CY;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_A_XOR;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_B;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_B1;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_B2;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_B3;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_B4;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_B5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_B6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_BO5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_BO6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_B_CY;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_B_XOR;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_C;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_C1;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_C2;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_C3;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_C4;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_C5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_C6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_CO5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_CO6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_C_CY;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_C_XOR;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_D;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_D1;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_D2;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_D3;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_D4;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_D5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_D6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_DO5;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_DO6;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_D_CY;
  wire [0:0] CLBLM_L_X78Y117_SLICE_X121Y117_D_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_AO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_A_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_BO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_B_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_CO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_C_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_DO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_DO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X120Y119_D_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_AO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_AO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_A_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_BO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_BO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_B_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_CO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_CO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_C_XOR;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D1;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D2;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D3;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D4;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_DO5;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_DO6;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D_CY;
  wire [0:0] CLBLM_L_X78Y119_SLICE_X121Y119_D_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_AO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_A_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_BO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_B_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_CO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_C_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_DO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_DO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X120Y120_D_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_AO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_AO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_A_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_BO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_BO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_B_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_CO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_CO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_C_XOR;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D1;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D2;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D3;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D4;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_DO5;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_DO6;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D_CY;
  wire [0:0] CLBLM_L_X78Y120_SLICE_X121Y120_D_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_AO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_A_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_BO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_BO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_B_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_CO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_CO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_C_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_DO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_DO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X120Y121_D_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_AO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_AO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_A_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_BO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_BO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_B_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_CO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_CO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_C_XOR;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D1;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D2;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D3;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D4;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_DO5;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_DO6;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D_CY;
  wire [0:0] CLBLM_L_X78Y121_SLICE_X121Y121_D_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_AO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_A_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_BO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_B_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_CO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_CO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_C_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_DO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_DO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X120Y122_D_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_AO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_AO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_A_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_BO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_BO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_B_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_CO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_CO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_C_XOR;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D1;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D2;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D3;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D4;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_DO5;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_DO6;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D_CY;
  wire [0:0] CLBLM_L_X78Y122_SLICE_X121Y122_D_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_AO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_A_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_BO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_B_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_CO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_C_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_DO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X120Y123_D_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_AO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_AO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_A_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_BO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_BO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_B_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_CO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_C_XOR;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D1;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D2;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D3;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D4;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_DO5;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_DO6;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D_CY;
  wire [0:0] CLBLM_L_X78Y123_SLICE_X121Y123_D_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_AO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_A_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_BO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_B_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_CO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_CO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_C_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_DO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_DO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X120Y124_D_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_AO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_AO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_A_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_BO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_BO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_B_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_CO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_CO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_C_XOR;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D1;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D2;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D3;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D4;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_DO5;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_DO6;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D_CY;
  wire [0:0] CLBLM_L_X78Y124_SLICE_X121Y124_D_XOR;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_A;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_A1;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_A2;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_A3;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_A4;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_A5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_A6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_AO5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_A_CY;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_A_XOR;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_B;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_B1;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_B2;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_B3;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_B4;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_B5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_B6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_BO5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_B_CY;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_B_XOR;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_C;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_C1;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_C2;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_C3;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_C4;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_C5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_C6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_CO5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_CO6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_C_CY;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_C_XOR;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_D;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_D1;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_D2;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_D3;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_D4;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_D5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_D6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_DO5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_DO6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_D_CY;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X120Y126_D_XOR;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_A;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_A1;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_A2;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_A3;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_A4;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_A5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_A6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_AO5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_AO6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_A_CY;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_A_XOR;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_B;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_B1;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_B2;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_B3;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_B4;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_B5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_B6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_BO5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_BO6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_B_CY;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_B_XOR;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_C;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_C1;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_C2;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_C3;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_C4;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_C5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_C6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_CO5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_CO6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_C_CY;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_C_XOR;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_D;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_D1;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_D2;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_D3;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_D4;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_D5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_D6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_DO5;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_DO6;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_D_CY;
  wire [0:0] CLBLM_L_X78Y126_SLICE_X121Y126_D_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_AO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_A_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_BO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_BO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_B_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_CO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_CO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_C_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_DO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_DO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X120Y129_D_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_AO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_AO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_A_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_BO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_BO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_B_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_CO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_CO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_C_XOR;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D1;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D2;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D3;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D4;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_DO5;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_DO6;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D_CY;
  wire [0:0] CLBLM_L_X78Y129_SLICE_X121Y129_D_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_AO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_A_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_BO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_BO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_B_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_CO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_CO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_C_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_DO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_DO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X154Y131_D_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_AO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_AO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_A_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_BO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_BO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_B_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_CO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_CO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_C_XOR;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D1;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D2;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D3;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D4;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_DO5;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_DO6;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D_CY;
  wire [0:0] CLBLM_L_X98Y131_SLICE_X155Y131_D_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_AO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_A_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_BO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_BO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_B_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_CO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_CO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_C_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_DO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_DO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X154Y132_D_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_AO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_AO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_A_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_BO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_BO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_B_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_CO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_CO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_C_XOR;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D1;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D2;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D3;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D4;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_DO5;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_DO6;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D_CY;
  wire [0:0] CLBLM_L_X98Y132_SLICE_X155Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AX;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CLK;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AMUX;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_XOR;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_A;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_A1;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_A2;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_A3;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_A4;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_A5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_A6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_AO5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_A_CY;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_A_XOR;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_B;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_B1;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_B2;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_B3;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_B4;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_B5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_B6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_BO5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_BO6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_B_CY;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_B_XOR;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_C;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_C1;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_C2;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_C3;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_C4;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_C5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_C6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_CO5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_CO6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_C_CY;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_C_XOR;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_D;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_D1;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_D2;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_D3;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_D4;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_D5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_D6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_DO5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_DO6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_D_CY;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X74Y116_D_XOR;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_A;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_A1;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_A2;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_A3;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_A4;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_A5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_A6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_AO5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_AO6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_A_CY;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_A_XOR;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_B;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_B1;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_B2;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_B3;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_B4;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_B5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_B6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_BO5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_BO6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_B_CY;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_B_XOR;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_C;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_C1;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_C2;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_C3;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_C4;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_C5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_C6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_CO5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_CO6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_C_CY;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_C_XOR;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_D;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_D1;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_D2;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_D3;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_D4;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_D5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_D6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_DO5;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_DO6;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_D_CY;
  wire [0:0] CLBLM_R_X49Y116_SLICE_X75Y116_D_XOR;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_A;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_A1;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_A2;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_A3;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_A4;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_A5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_A6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_AO5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_AO6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_AQ;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_AX;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_A_CY;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_A_XOR;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_B;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_B1;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_B2;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_B3;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_B4;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_B5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_B6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_BO5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_BO6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_B_CY;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_B_XOR;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_C;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_C1;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_C2;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_C3;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_C4;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_C5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_C6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_CLK;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_CO5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_CO6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_C_CY;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_C_XOR;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_D;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_D1;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_D2;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_D3;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_D4;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_D5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_D6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_DO5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_DO6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_D_CY;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X88Y117_D_XOR;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_A;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_A1;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_A2;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_A3;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_A4;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_A5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_A6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_AO5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_AO6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_A_CY;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_A_XOR;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_B;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_B1;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_B2;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_B3;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_B4;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_B5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_B6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_BO5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_BO6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_B_CY;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_B_XOR;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_C;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_C1;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_C2;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_C3;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_C4;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_C5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_C6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_CO5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_CO6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_C_CY;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_C_XOR;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_D;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_D1;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_D2;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_D3;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_D4;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_D5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_D6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_DO5;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_DO6;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_D_CY;
  wire [0:0] CLBLM_R_X59Y117_SLICE_X89Y117_D_XOR;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_A;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_A1;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_A2;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_A3;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_A4;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_A5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_A6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_AO5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_AO6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_AQ;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_AX;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_A_CY;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_A_XOR;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_B;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_B1;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_B2;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_B3;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_B4;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_B5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_B6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_BO5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_BO6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_B_CY;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_B_XOR;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_C;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_C1;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_C2;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_C3;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_C4;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_C5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_C6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_CLK;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_CO5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_CO6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_C_CY;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_C_XOR;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_D;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_D1;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_D2;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_D3;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_D4;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_D5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_D6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_DO5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_DO6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_D_CY;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X88Y118_D_XOR;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_A;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_A1;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_A2;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_A3;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_A4;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_A5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_A6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_AO5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_AO6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_A_CY;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_A_XOR;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_B;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_B1;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_B2;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_B3;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_B4;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_B5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_B6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_BO5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_BO6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_B_CY;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_B_XOR;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_C;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_C1;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_C2;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_C3;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_C4;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_C5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_C6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_CO5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_CO6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_C_CY;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_C_XOR;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_D;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_D1;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_D2;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_D3;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_D4;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_D5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_D6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_DO5;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_DO6;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_D_CY;
  wire [0:0] CLBLM_R_X59Y118_SLICE_X89Y118_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_I;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_I;
  wire [0:0] LIOB33_SING_X0Y200_IOB_X0Y200_I;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_SING_X0Y99_IOB_X0Y99_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_I;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_I;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_I;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_I;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_I;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_I;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_I;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_I;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_I;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_I;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_I;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_I;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_I;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_I;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_I;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_I;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_I;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_I;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_I;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_I;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_I;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_I;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_I;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_I;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_I;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y201_I;
  wire [0:0] LIOB33_X0Y201_IOB_X0Y202_I;
  wire [0:0] LIOB33_X0Y203_IOB_X0Y203_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y81_I;
  wire [0:0] LIOB33_X0Y81_IOB_X0Y82_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y83_I;
  wire [0:0] LIOB33_X0Y83_IOB_X0Y84_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y85_I;
  wire [0:0] LIOB33_X0Y85_IOB_X0Y86_O;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y87_O;
  wire [0:0] LIOB33_X0Y87_IOB_X0Y88_O;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y89_O;
  wire [0:0] LIOB33_X0Y89_IOB_X0Y90_O;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y91_O;
  wire [0:0] LIOB33_X0Y91_IOB_X0Y92_O;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y93_O;
  wire [0:0] LIOB33_X0Y93_IOB_X0Y94_O;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y95_O;
  wire [0:0] LIOB33_X0Y95_IOB_X0Y96_O;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y97_O;
  wire [0:0] LIOB33_X0Y97_IOB_X0Y98_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_D;
  wire [0:0] LIOI3_SING_X0Y150_ILOGIC_X0Y150_O;
  wire [0:0] LIOI3_SING_X0Y199_ILOGIC_X0Y199_D;
  wire [0:0] LIOI3_SING_X0Y199_ILOGIC_X0Y199_O;
  wire [0:0] LIOI3_SING_X0Y200_ILOGIC_X0Y200_D;
  wire [0:0] LIOI3_SING_X0Y200_ILOGIC_X0Y200_O;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_D1;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_OQ;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_T1;
  wire [0:0] LIOI3_SING_X0Y99_OLOGIC_X0Y99_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y151_O;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_D;
  wire [0:0] LIOI3_X0Y151_ILOGIC_X0Y152_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y153_O;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_D;
  wire [0:0] LIOI3_X0Y153_ILOGIC_X0Y154_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y155_O;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_D;
  wire [0:0] LIOI3_X0Y155_ILOGIC_X0Y156_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y159_O;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_D;
  wire [0:0] LIOI3_X0Y159_ILOGIC_X0Y160_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y161_O;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_D;
  wire [0:0] LIOI3_X0Y161_ILOGIC_X0Y162_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y165_O;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_D;
  wire [0:0] LIOI3_X0Y165_ILOGIC_X0Y166_O;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y167_D;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y167_O;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_D;
  wire [0:0] LIOI3_X0Y167_ILOGIC_X0Y168_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y171_O;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_D;
  wire [0:0] LIOI3_X0Y171_ILOGIC_X0Y172_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y173_O;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_D;
  wire [0:0] LIOI3_X0Y173_ILOGIC_X0Y174_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y175_O;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_D;
  wire [0:0] LIOI3_X0Y175_ILOGIC_X0Y176_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y177_O;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_D;
  wire [0:0] LIOI3_X0Y177_ILOGIC_X0Y178_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y179_O;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_D;
  wire [0:0] LIOI3_X0Y179_ILOGIC_X0Y180_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y183_O;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_D;
  wire [0:0] LIOI3_X0Y183_ILOGIC_X0Y184_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y185_O;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_D;
  wire [0:0] LIOI3_X0Y185_ILOGIC_X0Y186_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y189_O;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_D;
  wire [0:0] LIOI3_X0Y189_ILOGIC_X0Y190_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y191_O;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_D;
  wire [0:0] LIOI3_X0Y191_ILOGIC_X0Y192_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y195_O;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_D;
  wire [0:0] LIOI3_X0Y195_ILOGIC_X0Y196_O;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_D;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y197_O;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y198_D;
  wire [0:0] LIOI3_X0Y197_ILOGIC_X0Y198_O;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y201_D;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y201_O;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y202_D;
  wire [0:0] LIOI3_X0Y201_ILOGIC_X0Y202_O;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y203_D;
  wire [0:0] LIOI3_X0Y203_ILOGIC_X0Y203_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y80_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y83_O;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_D;
  wire [0:0] LIOI3_X0Y83_ILOGIC_X0Y84_O;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_D;
  wire [0:0] LIOI3_X0Y85_ILOGIC_X0Y85_O;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_D1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_OQ;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_T1;
  wire [0:0] LIOI3_X0Y85_OLOGIC_X0Y86_TQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_D1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_OQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_T1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y89_TQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_D1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_OQ;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_T1;
  wire [0:0] LIOI3_X0Y89_OLOGIC_X0Y90_TQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_D1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_OQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_T1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y91_TQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_D1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_OQ;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_T1;
  wire [0:0] LIOI3_X0Y91_OLOGIC_X0Y92_TQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_D1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_OQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_T1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y95_TQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_D1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_OQ;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_T1;
  wire [0:0] LIOI3_X0Y95_OLOGIC_X0Y96_TQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_D1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_OQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_T1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y97_TQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_D1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_OQ;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_T1;
  wire [0:0] LIOI3_X0Y97_OLOGIC_X0Y98_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_I;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_I;
  wire [0:0] RIOB33_SING_X105Y50_IOB_X1Y50_I;
  wire [0:0] RIOB33_SING_X105Y99_IOB_X1Y99_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_I;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_I;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_I;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_I;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_I;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_I;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_I;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_I;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_I;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_I;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_I;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_I;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_I;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_I;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_I;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_I;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_I;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_I;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_I;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_I;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_I;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_I;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_I;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_I;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_I;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_I;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_I;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_I;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_I;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_I;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_I;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_I;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_I;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_I;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_I;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_I;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_I;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_I;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_I;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_I;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_I;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_I;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_I;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_I;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_I;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_I;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_I;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y51_I;
  wire [0:0] RIOB33_X105Y51_IOB_X1Y52_I;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y53_I;
  wire [0:0] RIOB33_X105Y53_IOB_X1Y54_I;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y55_I;
  wire [0:0] RIOB33_X105Y55_IOB_X1Y56_I;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y57_I;
  wire [0:0] RIOB33_X105Y57_IOB_X1Y58_I;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y59_I;
  wire [0:0] RIOB33_X105Y59_IOB_X1Y60_I;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y61_I;
  wire [0:0] RIOB33_X105Y61_IOB_X1Y62_I;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y63_I;
  wire [0:0] RIOB33_X105Y63_IOB_X1Y64_I;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y65_I;
  wire [0:0] RIOB33_X105Y65_IOB_X1Y66_I;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y67_I;
  wire [0:0] RIOB33_X105Y67_IOB_X1Y68_I;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y69_I;
  wire [0:0] RIOB33_X105Y69_IOB_X1Y70_I;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y71_I;
  wire [0:0] RIOB33_X105Y71_IOB_X1Y72_I;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y73_I;
  wire [0:0] RIOB33_X105Y73_IOB_X1Y74_I;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y75_I;
  wire [0:0] RIOB33_X105Y75_IOB_X1Y76_I;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y77_I;
  wire [0:0] RIOB33_X105Y77_IOB_X1Y78_I;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y79_I;
  wire [0:0] RIOB33_X105Y79_IOB_X1Y80_I;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y81_I;
  wire [0:0] RIOB33_X105Y81_IOB_X1Y82_I;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y83_I;
  wire [0:0] RIOB33_X105Y83_IOB_X1Y84_I;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y85_I;
  wire [0:0] RIOB33_X105Y85_IOB_X1Y86_I;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y87_I;
  wire [0:0] RIOB33_X105Y87_IOB_X1Y88_I;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y89_I;
  wire [0:0] RIOB33_X105Y89_IOB_X1Y90_I;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y91_I;
  wire [0:0] RIOB33_X105Y91_IOB_X1Y92_I;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y93_I;
  wire [0:0] RIOB33_X105Y93_IOB_X1Y94_I;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y95_I;
  wire [0:0] RIOB33_X105Y95_IOB_X1Y96_I;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y97_I;
  wire [0:0] RIOB33_X105Y97_IOB_X1Y98_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_ILOGIC_X1Y150_D;
  wire [0:0] RIOI3_SING_X105Y150_ILOGIC_X1Y150_O;
  wire [0:0] RIOI3_SING_X105Y199_ILOGIC_X1Y199_D;
  wire [0:0] RIOI3_SING_X105Y199_ILOGIC_X1Y199_O;
  wire [0:0] RIOI3_SING_X105Y50_ILOGIC_X1Y50_D;
  wire [0:0] RIOI3_SING_X105Y50_ILOGIC_X1Y50_O;
  wire [0:0] RIOI3_SING_X105Y99_ILOGIC_X1Y99_D;
  wire [0:0] RIOI3_SING_X105Y99_ILOGIC_X1Y99_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y181_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y181_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y182_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y182_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y193_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y193_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y194_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y194_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y57_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y57_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y58_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y58_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_ILOGIC_X1Y69_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_ILOGIC_X1Y69_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_ILOGIC_X1Y70_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y69_ILOGIC_X1Y70_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_ILOGIC_X1Y81_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_ILOGIC_X1Y81_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_ILOGIC_X1Y82_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y81_ILOGIC_X1Y82_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_ILOGIC_X1Y93_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_ILOGIC_X1Y93_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_ILOGIC_X1Y94_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y93_ILOGIC_X1Y94_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y164_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y164_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y187_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y187_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y188_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y188_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_ILOGIC_X1Y63_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_ILOGIC_X1Y63_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_ILOGIC_X1Y64_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y63_ILOGIC_X1Y64_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_ILOGIC_X1Y87_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_ILOGIC_X1Y87_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_ILOGIC_X1Y88_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y87_ILOGIC_X1Y88_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y151_D;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y151_O;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y152_D;
  wire [0:0] RIOI3_X105Y151_ILOGIC_X1Y152_O;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y153_D;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y153_O;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y154_D;
  wire [0:0] RIOI3_X105Y153_ILOGIC_X1Y154_O;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y155_D;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y155_O;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y156_D;
  wire [0:0] RIOI3_X105Y155_ILOGIC_X1Y156_O;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y159_D;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y159_O;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y160_D;
  wire [0:0] RIOI3_X105Y159_ILOGIC_X1Y160_O;
  wire [0:0] RIOI3_X105Y161_ILOGIC_X1Y161_D;
  wire [0:0] RIOI3_X105Y161_ILOGIC_X1Y161_O;
  wire [0:0] RIOI3_X105Y161_ILOGIC_X1Y162_D;
  wire [0:0] RIOI3_X105Y161_ILOGIC_X1Y162_O;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y165_D;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y165_O;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y166_D;
  wire [0:0] RIOI3_X105Y165_ILOGIC_X1Y166_O;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y167_D;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y167_O;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y168_D;
  wire [0:0] RIOI3_X105Y167_ILOGIC_X1Y168_O;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y171_D;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y171_O;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y172_D;
  wire [0:0] RIOI3_X105Y171_ILOGIC_X1Y172_O;
  wire [0:0] RIOI3_X105Y173_ILOGIC_X1Y173_D;
  wire [0:0] RIOI3_X105Y173_ILOGIC_X1Y173_O;
  wire [0:0] RIOI3_X105Y173_ILOGIC_X1Y174_D;
  wire [0:0] RIOI3_X105Y173_ILOGIC_X1Y174_O;
  wire [0:0] RIOI3_X105Y175_ILOGIC_X1Y175_D;
  wire [0:0] RIOI3_X105Y175_ILOGIC_X1Y175_O;
  wire [0:0] RIOI3_X105Y175_ILOGIC_X1Y176_D;
  wire [0:0] RIOI3_X105Y175_ILOGIC_X1Y176_O;
  wire [0:0] RIOI3_X105Y177_ILOGIC_X1Y177_D;
  wire [0:0] RIOI3_X105Y177_ILOGIC_X1Y177_O;
  wire [0:0] RIOI3_X105Y177_ILOGIC_X1Y178_D;
  wire [0:0] RIOI3_X105Y177_ILOGIC_X1Y178_O;
  wire [0:0] RIOI3_X105Y179_ILOGIC_X1Y179_D;
  wire [0:0] RIOI3_X105Y179_ILOGIC_X1Y179_O;
  wire [0:0] RIOI3_X105Y179_ILOGIC_X1Y180_D;
  wire [0:0] RIOI3_X105Y179_ILOGIC_X1Y180_O;
  wire [0:0] RIOI3_X105Y183_ILOGIC_X1Y183_D;
  wire [0:0] RIOI3_X105Y183_ILOGIC_X1Y183_O;
  wire [0:0] RIOI3_X105Y183_ILOGIC_X1Y184_D;
  wire [0:0] RIOI3_X105Y183_ILOGIC_X1Y184_O;
  wire [0:0] RIOI3_X105Y185_ILOGIC_X1Y185_D;
  wire [0:0] RIOI3_X105Y185_ILOGIC_X1Y185_O;
  wire [0:0] RIOI3_X105Y185_ILOGIC_X1Y186_D;
  wire [0:0] RIOI3_X105Y185_ILOGIC_X1Y186_O;
  wire [0:0] RIOI3_X105Y189_ILOGIC_X1Y189_D;
  wire [0:0] RIOI3_X105Y189_ILOGIC_X1Y189_O;
  wire [0:0] RIOI3_X105Y189_ILOGIC_X1Y190_D;
  wire [0:0] RIOI3_X105Y189_ILOGIC_X1Y190_O;
  wire [0:0] RIOI3_X105Y191_ILOGIC_X1Y191_D;
  wire [0:0] RIOI3_X105Y191_ILOGIC_X1Y191_O;
  wire [0:0] RIOI3_X105Y191_ILOGIC_X1Y192_D;
  wire [0:0] RIOI3_X105Y191_ILOGIC_X1Y192_O;
  wire [0:0] RIOI3_X105Y195_ILOGIC_X1Y195_D;
  wire [0:0] RIOI3_X105Y195_ILOGIC_X1Y195_O;
  wire [0:0] RIOI3_X105Y195_ILOGIC_X1Y196_D;
  wire [0:0] RIOI3_X105Y195_ILOGIC_X1Y196_O;
  wire [0:0] RIOI3_X105Y197_ILOGIC_X1Y197_D;
  wire [0:0] RIOI3_X105Y197_ILOGIC_X1Y197_O;
  wire [0:0] RIOI3_X105Y197_ILOGIC_X1Y198_D;
  wire [0:0] RIOI3_X105Y197_ILOGIC_X1Y198_O;
  wire [0:0] RIOI3_X105Y51_ILOGIC_X1Y51_D;
  wire [0:0] RIOI3_X105Y51_ILOGIC_X1Y51_O;
  wire [0:0] RIOI3_X105Y51_ILOGIC_X1Y52_D;
  wire [0:0] RIOI3_X105Y51_ILOGIC_X1Y52_O;
  wire [0:0] RIOI3_X105Y53_ILOGIC_X1Y53_D;
  wire [0:0] RIOI3_X105Y53_ILOGIC_X1Y53_O;
  wire [0:0] RIOI3_X105Y53_ILOGIC_X1Y54_D;
  wire [0:0] RIOI3_X105Y53_ILOGIC_X1Y54_O;
  wire [0:0] RIOI3_X105Y55_ILOGIC_X1Y55_D;
  wire [0:0] RIOI3_X105Y55_ILOGIC_X1Y55_O;
  wire [0:0] RIOI3_X105Y55_ILOGIC_X1Y56_D;
  wire [0:0] RIOI3_X105Y55_ILOGIC_X1Y56_O;
  wire [0:0] RIOI3_X105Y59_ILOGIC_X1Y59_D;
  wire [0:0] RIOI3_X105Y59_ILOGIC_X1Y59_O;
  wire [0:0] RIOI3_X105Y59_ILOGIC_X1Y60_D;
  wire [0:0] RIOI3_X105Y59_ILOGIC_X1Y60_O;
  wire [0:0] RIOI3_X105Y61_ILOGIC_X1Y61_D;
  wire [0:0] RIOI3_X105Y61_ILOGIC_X1Y61_O;
  wire [0:0] RIOI3_X105Y61_ILOGIC_X1Y62_D;
  wire [0:0] RIOI3_X105Y61_ILOGIC_X1Y62_O;
  wire [0:0] RIOI3_X105Y65_ILOGIC_X1Y65_D;
  wire [0:0] RIOI3_X105Y65_ILOGIC_X1Y65_O;
  wire [0:0] RIOI3_X105Y65_ILOGIC_X1Y66_D;
  wire [0:0] RIOI3_X105Y65_ILOGIC_X1Y66_O;
  wire [0:0] RIOI3_X105Y67_ILOGIC_X1Y67_D;
  wire [0:0] RIOI3_X105Y67_ILOGIC_X1Y67_O;
  wire [0:0] RIOI3_X105Y67_ILOGIC_X1Y68_D;
  wire [0:0] RIOI3_X105Y67_ILOGIC_X1Y68_O;
  wire [0:0] RIOI3_X105Y71_ILOGIC_X1Y71_D;
  wire [0:0] RIOI3_X105Y71_ILOGIC_X1Y71_O;
  wire [0:0] RIOI3_X105Y71_ILOGIC_X1Y72_D;
  wire [0:0] RIOI3_X105Y71_ILOGIC_X1Y72_O;
  wire [0:0] RIOI3_X105Y73_ILOGIC_X1Y73_D;
  wire [0:0] RIOI3_X105Y73_ILOGIC_X1Y73_O;
  wire [0:0] RIOI3_X105Y73_ILOGIC_X1Y74_D;
  wire [0:0] RIOI3_X105Y73_ILOGIC_X1Y74_O;
  wire [0:0] RIOI3_X105Y75_ILOGIC_X1Y75_D;
  wire [0:0] RIOI3_X105Y75_ILOGIC_X1Y75_O;
  wire [0:0] RIOI3_X105Y75_ILOGIC_X1Y76_D;
  wire [0:0] RIOI3_X105Y75_ILOGIC_X1Y76_O;
  wire [0:0] RIOI3_X105Y77_ILOGIC_X1Y77_D;
  wire [0:0] RIOI3_X105Y77_ILOGIC_X1Y77_O;
  wire [0:0] RIOI3_X105Y77_ILOGIC_X1Y78_D;
  wire [0:0] RIOI3_X105Y77_ILOGIC_X1Y78_O;
  wire [0:0] RIOI3_X105Y79_ILOGIC_X1Y79_D;
  wire [0:0] RIOI3_X105Y79_ILOGIC_X1Y79_O;
  wire [0:0] RIOI3_X105Y79_ILOGIC_X1Y80_D;
  wire [0:0] RIOI3_X105Y79_ILOGIC_X1Y80_O;
  wire [0:0] RIOI3_X105Y83_ILOGIC_X1Y83_D;
  wire [0:0] RIOI3_X105Y83_ILOGIC_X1Y83_O;
  wire [0:0] RIOI3_X105Y83_ILOGIC_X1Y84_D;
  wire [0:0] RIOI3_X105Y83_ILOGIC_X1Y84_O;
  wire [0:0] RIOI3_X105Y85_ILOGIC_X1Y85_D;
  wire [0:0] RIOI3_X105Y85_ILOGIC_X1Y85_O;
  wire [0:0] RIOI3_X105Y85_ILOGIC_X1Y86_D;
  wire [0:0] RIOI3_X105Y85_ILOGIC_X1Y86_O;
  wire [0:0] RIOI3_X105Y89_ILOGIC_X1Y89_D;
  wire [0:0] RIOI3_X105Y89_ILOGIC_X1Y89_O;
  wire [0:0] RIOI3_X105Y89_ILOGIC_X1Y90_D;
  wire [0:0] RIOI3_X105Y89_ILOGIC_X1Y90_O;
  wire [0:0] RIOI3_X105Y91_ILOGIC_X1Y91_D;
  wire [0:0] RIOI3_X105Y91_ILOGIC_X1Y91_O;
  wire [0:0] RIOI3_X105Y91_ILOGIC_X1Y92_D;
  wire [0:0] RIOI3_X105Y91_ILOGIC_X1Y92_O;
  wire [0:0] RIOI3_X105Y95_ILOGIC_X1Y95_D;
  wire [0:0] RIOI3_X105Y95_ILOGIC_X1Y95_O;
  wire [0:0] RIOI3_X105Y95_ILOGIC_X1Y96_D;
  wire [0:0] RIOI3_X105Y95_ILOGIC_X1Y96_O;
  wire [0:0] RIOI3_X105Y97_ILOGIC_X1Y97_D;
  wire [0:0] RIOI3_X105Y97_ILOGIC_X1Y97_O;
  wire [0:0] RIOI3_X105Y97_ILOGIC_X1Y98_D;
  wire [0:0] RIOI3_X105Y97_ILOGIC_X1Y98_O;


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.Q(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X0Y105_CO6),
.Q(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.Q(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f3eec022)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_DLUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I5(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c393c6c)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(CLBLL_R_X71Y116_SLICE_X107Y116_AO6),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.I3(LIOB33_X0Y81_IOB_X0Y82_I),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y80_I),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc0300fece3202)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_BLUT (
.I0(LIOB33_X0Y51_IOB_X0Y51_I),
.I1(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001fffdfffe0002)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_ALUT (
.I0(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(LIOB33_X0Y79_IOB_X0Y80_I),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I5(CLBLL_R_X71Y120_SLICE_X107Y120_CO6),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050fbea5140)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I4(LIOB33_X0Y53_IOB_X0Y54_I),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fb51fa50ea40)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I3(LIOB33_X0Y51_IOB_X0Y52_I),
.I4(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y118_SLICE_X0Y118_CO6),
.Q(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.Q(CLBLL_L_X2Y118_SLICE_X0Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfcfa0c0a)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_CLUT (
.I0(CLBLL_L_X2Y118_SLICE_X0Y118_BQ),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I2(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e4f0e4f0ddf088)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLL_L_X2Y118_SLICE_X0Y118_BQ),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(LIOB33_X0Y75_IOB_X0Y76_I),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e1ff0f0f1e0)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(CLBLL_L_X2Y118_SLICE_X0Y118_AQ),
.I3(CLBLL_L_X2Y118_SLICE_X0Y118_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_R_X71Y118_SLICE_X106Y118_AO6),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.Q(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.Q(CLBLL_L_X2Y119_SLICE_X0Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444efea4540)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I1(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.I2(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_BQ),
.I4(LIOB33_X0Y57_IOB_X0Y57_I),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e4ddf0f0e488)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(CLBLL_L_X2Y119_SLICE_X0Y119_BQ),
.I2(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I5(LIOB33_X0Y55_IOB_X0Y56_I),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e1ff0f0f1e0)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLL_L_X2Y119_SLICE_X0Y119_AQ),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y80_I),
.I5(CLBLM_L_X68Y119_SLICE_X103Y119_BO6),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.Q(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.Q(CLBLL_L_X2Y119_SLICE_X1Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0f3e2c0e2)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_BQ),
.I1(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I2(LIOB33_X0Y71_IOB_X0Y71_I),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e4ddf0f0e488)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_BQ),
.I2(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I5(LIOB33_X0Y69_IOB_X0Y70_I),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h666666666666636c)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I1(CLBLM_L_X68Y119_SLICE_X103Y119_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y80_I),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.Q(CLBLL_L_X2Y120_SLICE_X0Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.Q(CLBLL_L_X2Y120_SLICE_X0Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888ddd88d88)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I1(LIOB33_X0Y69_IOB_X0Y69_I),
.I2(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000cccaccca)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(CLBLL_L_X2Y120_SLICE_X0Y120_BQ),
.I1(CLBLL_L_X2Y120_SLICE_X0Y120_AQ),
.I2(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffca000c00ca)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLL_L_X2Y120_SLICE_X0Y120_BQ),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(CLBLL_L_X2Y120_SLICE_X0Y120_AQ),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a596a)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(CLBLL_R_X71Y119_SLICE_X106Y119_DO6),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(CLBLL_L_X2Y120_SLICE_X0Y120_AQ),
.I3(CLBLL_L_X2Y120_SLICE_X0Y120_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(LIOB33_X0Y79_IOB_X0Y80_I),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.Q(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3e2c0d1c0c0)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_DLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I1(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I2(LIOB33_X0Y73_IOB_X0Y73_I),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(CLBLL_L_X2Y123_SLICE_X0Y123_DQ),
.I5(CLBLL_L_X2Y123_SLICE_X0Y123_BQ),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeedec13120100)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_CLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(LIOB33_X0Y71_IOB_X0Y72_I),
.I4(CLBLL_L_X2Y123_SLICE_X0Y123_DQ),
.I5(CLBLL_L_X2Y123_SLICE_X0Y123_BQ),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fec23e02)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I5(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001fefffffe0100)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(LIOB33_X0Y79_IOB_X0Y80_I),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I5(CLBLM_L_X68Y119_SLICE_X103Y119_AO6),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y123_SLICE_X0Y123_CO6),
.Q(CLBLL_L_X2Y123_SLICE_X0Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y121_SLICE_X0Y121_DO6),
.Q(CLBLL_L_X2Y123_SLICE_X0Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y123_SLICE_X0Y123_AO6),
.Q(CLBLL_L_X2Y123_SLICE_X0Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_AO6),
.Q(CLBLL_L_X2Y123_SLICE_X0Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff11ee00)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_DLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I2(LIOB33_X0Y75_IOB_X0Y75_I),
.I3(CLBLL_L_X2Y124_SLICE_X0Y124_AQ),
.I4(CLBLL_L_X2Y124_SLICE_X0Y124_CQ),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0e4f0e4)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_CLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I1(CLBLL_L_X2Y123_SLICE_X0Y123_CQ),
.I2(CLBLL_L_X2Y123_SLICE_X0Y123_AQ),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(LIOB33_X0Y67_IOB_X0Y67_I),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f3c0ee22)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_BLUT (
.I0(LIOB33_X0Y65_IOB_X0Y66_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(CLBLL_L_X2Y123_SLICE_X0Y123_AQ),
.I3(CLBLL_L_X2Y123_SLICE_X0Y123_CQ),
.I4(LIOB33_X0Y83_IOB_X0Y83_I),
.I5(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e1ff0f0f1e0)
  ) CLBLL_L_X2Y123_SLICE_X0Y123_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLL_L_X2Y123_SLICE_X0Y123_AQ),
.I3(CLBLL_L_X2Y123_SLICE_X0Y123_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLL_R_X71Y120_SLICE_X107Y120_BO6),
.O5(CLBLL_L_X2Y123_SLICE_X0Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X0Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_DO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_CO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccfccfaccc0cc0a)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_BLUT (
.I0(LIOB33_X0Y73_IOB_X0Y74_I),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_AQ),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(CLBLL_L_X2Y124_SLICE_X0Y124_CQ),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_BO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00fe32ce02)
  ) CLBLL_L_X2Y123_SLICE_X1Y123_ALUT (
.I0(CLBLL_L_X2Y124_SLICE_X1Y124_DQ),
.I1(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I2(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I3(LIOB33_X0Y61_IOB_X0Y61_I),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.O5(CLBLL_L_X2Y123_SLICE_X1Y123_AO5),
.O6(CLBLL_L_X2Y123_SLICE_X1Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y123_SLICE_X0Y123_DO6),
.Q(CLBLL_L_X2Y124_SLICE_X0Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y124_SLICE_X0Y124_CO6),
.Q(CLBLL_L_X2Y124_SLICE_X0Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.Q(CLBLL_L_X2Y124_SLICE_X0Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y124_SLICE_X0Y124_AO6),
.Q(CLBLL_L_X2Y124_SLICE_X0Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0f3e2d1c0)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_DLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I1(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I2(LIOB33_X0Y65_IOB_X0Y65_I),
.I3(CLBLL_L_X2Y124_SLICE_X1Y124_CQ),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_BQ),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_DO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeefc22222230)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_CLUT (
.I0(CLBLL_L_X2Y124_SLICE_X0Y124_BQ),
.I1(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I2(CLBLL_L_X2Y124_SLICE_X0Y124_DQ),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I5(LIOB33_X0Y63_IOB_X0Y63_I),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_CO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe030efcf20002)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(CLBLL_L_X2Y124_SLICE_X0Y124_BQ),
.I5(CLBLL_L_X2Y124_SLICE_X0Y124_DQ),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_BO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333237cccccdc8)
  ) CLBLL_L_X2Y124_SLICE_X0Y124_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(CLBLL_L_X2Y124_SLICE_X0Y124_BQ),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(CLBLL_L_X2Y124_SLICE_X0Y124_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y80_I),
.I5(CLBLL_R_X71Y126_SLICE_X106Y126_AO6),
.O5(CLBLL_L_X2Y124_SLICE_X0Y124_AO5),
.O6(CLBLL_L_X2Y124_SLICE_X0Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.Q(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.Q(CLBLL_L_X2Y124_SLICE_X1Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y124_SLICE_X1Y124_CO6),
.Q(CLBLL_L_X2Y124_SLICE_X1Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y124_SLICE_X1Y124_AO6),
.Q(CLBLL_L_X2Y124_SLICE_X1Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0e4dde488)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_DLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLL_L_X2Y124_SLICE_X1Y124_CQ),
.I2(CLBLL_L_X2Y124_SLICE_X1Y124_BQ),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(LIOB33_X0Y63_IOB_X0Y64_I),
.I5(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_DO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c393c6c)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(CLBLL_R_X71Y126_SLICE_X106Y126_BO6),
.I2(CLBLL_L_X2Y124_SLICE_X1Y124_BQ),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(CLBLL_L_X2Y124_SLICE_X1Y124_DO6),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_CO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f0eef0c0f022)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_BLUT (
.I0(LIOB33_X0Y59_IOB_X0Y60_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(LIOB33_X0Y83_IOB_X0Y83_I),
.I5(CLBLL_L_X2Y124_SLICE_X1Y124_DQ),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_BO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a596a)
  ) CLBLL_L_X2Y124_SLICE_X1Y124_ALUT (
.I0(CLBLL_R_X71Y125_SLICE_X106Y125_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(CLBLL_L_X2Y124_SLICE_X1Y124_AQ),
.I3(CLBLL_L_X2Y124_SLICE_X1Y124_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_L_X2Y124_SLICE_X1Y124_AO5),
.O6(CLBLL_L_X2Y124_SLICE_X1Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaafff000f0)
  ) CLBLL_R_X71Y116_SLICE_X106Y116_DLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X71Y116_SLICE_X106Y116_DO5),
.O6(CLBLL_R_X71Y116_SLICE_X106Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0aaccaacc)
  ) CLBLL_R_X71Y116_SLICE_X106Y116_CLUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X71Y116_SLICE_X106Y116_CO5),
.O6(CLBLL_R_X71Y116_SLICE_X106Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bb88bb88)
  ) CLBLL_R_X71Y116_SLICE_X106Y116_BLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLL_R_X71Y116_SLICE_X106Y116_BO5),
.O6(CLBLL_R_X71Y116_SLICE_X106Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbfc308888fc30)
  ) CLBLL_R_X71Y116_SLICE_X106Y116_ALUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.O5(CLBLL_R_X71Y116_SLICE_X106Y116_AO5),
.O6(CLBLL_R_X71Y116_SLICE_X106Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y116_SLICE_X106Y116_MUXF7A (
.I0(CLBLL_R_X71Y116_SLICE_X106Y116_BO6),
.I1(CLBLL_R_X71Y116_SLICE_X106Y116_AO6),
.O(CLBLL_R_X71Y116_SLICE_X106Y116_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y116_SLICE_X106Y116_MUXF7B (
.I0(CLBLL_R_X71Y116_SLICE_X106Y116_DO6),
.I1(CLBLL_R_X71Y116_SLICE_X106Y116_CO6),
.O(CLBLL_R_X71Y116_SLICE_X106Y116_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X71Y116_SLICE_X106Y116_MUXF8 (
.I0(CLBLL_R_X71Y116_SLICE_X106Y116_F7BMUX_O),
.I1(CLBLL_R_X71Y116_SLICE_X106Y116_F7AMUX_O),
.O(CLBLL_R_X71Y116_SLICE_X106Y116_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5f2da2569199693)
  ) CLBLL_R_X71Y116_SLICE_X107Y116_DLUT (
.I0(CLBLL_R_X73Y115_SLICE_X110Y115_CO6),
.I1(CLBLM_L_X74Y116_SLICE_X113Y116_CO6),
.I2(CLBLM_L_X72Y119_SLICE_X108Y119_DO6),
.I3(CLBLM_L_X72Y119_SLICE_X108Y119_CO6),
.I4(CLBLL_R_X75Y116_SLICE_X114Y116_CO6),
.I5(CLBLM_L_X72Y116_SLICE_X108Y116_CO6),
.O5(CLBLL_R_X71Y116_SLICE_X107Y116_DO5),
.O6(CLBLL_R_X71Y116_SLICE_X107Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcb352d5a69866669)
  ) CLBLL_R_X71Y116_SLICE_X107Y116_CLUT (
.I0(CLBLL_R_X73Y115_SLICE_X110Y115_CO6),
.I1(CLBLM_L_X74Y116_SLICE_X113Y116_CO6),
.I2(CLBLM_L_X72Y116_SLICE_X108Y116_CO6),
.I3(CLBLM_L_X72Y119_SLICE_X108Y119_CO6),
.I4(CLBLL_R_X75Y116_SLICE_X114Y116_CO6),
.I5(CLBLM_L_X72Y119_SLICE_X108Y119_DO6),
.O5(CLBLL_R_X71Y116_SLICE_X107Y116_CO5),
.O6(CLBLL_R_X71Y116_SLICE_X107Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h635ce916589797a8)
  ) CLBLL_R_X71Y116_SLICE_X107Y116_BLUT (
.I0(CLBLM_L_X72Y116_SLICE_X108Y116_CO6),
.I1(CLBLM_L_X74Y116_SLICE_X113Y116_CO6),
.I2(CLBLM_L_X72Y119_SLICE_X108Y119_CO6),
.I3(CLBLM_L_X72Y119_SLICE_X108Y119_DO6),
.I4(CLBLL_R_X73Y115_SLICE_X110Y115_CO6),
.I5(CLBLL_R_X75Y116_SLICE_X114Y116_CO6),
.O5(CLBLL_R_X71Y116_SLICE_X107Y116_BO5),
.O6(CLBLL_R_X71Y116_SLICE_X107Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc636398d2ed29cd2)
  ) CLBLL_R_X71Y116_SLICE_X107Y116_ALUT (
.I0(CLBLM_L_X72Y116_SLICE_X108Y116_CO6),
.I1(CLBLM_L_X74Y116_SLICE_X113Y116_CO6),
.I2(CLBLM_L_X72Y119_SLICE_X108Y119_CO6),
.I3(CLBLM_L_X72Y119_SLICE_X108Y119_DO6),
.I4(CLBLL_R_X73Y115_SLICE_X110Y115_CO6),
.I5(CLBLL_R_X75Y116_SLICE_X114Y116_CO6),
.O5(CLBLL_R_X71Y116_SLICE_X107Y116_AO5),
.O6(CLBLL_R_X71Y116_SLICE_X107Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4ffaae4e45500)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_DLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.O5(CLBLL_R_X71Y117_SLICE_X106Y117_DO5),
.O6(CLBLL_R_X71Y117_SLICE_X106Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe4aae455e400e4)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_CLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.O5(CLBLL_R_X71Y117_SLICE_X106Y117_CO5),
.O6(CLBLL_R_X71Y117_SLICE_X106Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfa0cfafc0a0c0a)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_BLUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I5(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.O5(CLBLL_R_X71Y117_SLICE_X106Y117_BO5),
.O6(CLBLL_R_X71Y117_SLICE_X106Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffacf0ac0fac00ac)
  ) CLBLL_R_X71Y117_SLICE_X106Y117_ALUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I1(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.O5(CLBLL_R_X71Y117_SLICE_X106Y117_AO5),
.O6(CLBLL_R_X71Y117_SLICE_X106Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y117_SLICE_X106Y117_MUXF7A (
.I0(CLBLL_R_X71Y117_SLICE_X106Y117_BO6),
.I1(CLBLL_R_X71Y117_SLICE_X106Y117_AO6),
.O(CLBLL_R_X71Y117_SLICE_X106Y117_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y117_SLICE_X106Y117_MUXF7B (
.I0(CLBLL_R_X71Y117_SLICE_X106Y117_DO6),
.I1(CLBLL_R_X71Y117_SLICE_X106Y117_CO6),
.O(CLBLL_R_X71Y117_SLICE_X106Y117_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X107Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X107Y117_DO5),
.O6(CLBLL_R_X71Y117_SLICE_X107Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X107Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X107Y117_CO5),
.O6(CLBLL_R_X71Y117_SLICE_X107Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X107Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X107Y117_BO5),
.O6(CLBLL_R_X71Y117_SLICE_X107Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y117_SLICE_X107Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y117_SLICE_X107Y117_AO5),
.O6(CLBLL_R_X71Y117_SLICE_X107Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y118_SLICE_X106Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y118_SLICE_X106Y118_DO5),
.O6(CLBLL_R_X71Y118_SLICE_X106Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y118_SLICE_X106Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y118_SLICE_X106Y118_CO5),
.O6(CLBLL_R_X71Y118_SLICE_X106Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y118_SLICE_X106Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y118_SLICE_X106Y118_BO5),
.O6(CLBLL_R_X71Y118_SLICE_X106Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h703996e64f94e836)
  ) CLBLL_R_X71Y118_SLICE_X106Y118_ALUT (
.I0(CLBLM_L_X74Y117_SLICE_X113Y117_DO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_CO6),
.I2(CLBLM_L_X74Y117_SLICE_X113Y117_CO6),
.I3(CLBLL_R_X73Y116_SLICE_X110Y116_CO6),
.I4(CLBLM_L_X72Y116_SLICE_X108Y116_DO6),
.I5(CLBLL_R_X75Y120_SLICE_X115Y120_CO6),
.O5(CLBLL_R_X71Y118_SLICE_X106Y118_AO5),
.O6(CLBLL_R_X71Y118_SLICE_X106Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50dddd8888)
  ) CLBLL_R_X71Y118_SLICE_X107Y118_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I4(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLL_R_X71Y118_SLICE_X107Y118_DO5),
.O6(CLBLL_R_X71Y118_SLICE_X107Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef4aea45e540e04)
  ) CLBLL_R_X71Y118_SLICE_X107Y118_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I4(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.O5(CLBLL_R_X71Y118_SLICE_X107Y118_CO5),
.O6(CLBLL_R_X71Y118_SLICE_X107Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfceefc2230ee3022)
  ) CLBLL_R_X71Y118_SLICE_X107Y118_BLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.O5(CLBLL_R_X71Y118_SLICE_X107Y118_BO5),
.O6(CLBLL_R_X71Y118_SLICE_X107Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffac0facf0ac00ac)
  ) CLBLL_R_X71Y118_SLICE_X107Y118_ALUT (
.I0(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I5(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.O5(CLBLL_R_X71Y118_SLICE_X107Y118_AO5),
.O6(CLBLL_R_X71Y118_SLICE_X107Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y118_SLICE_X107Y118_MUXF7A (
.I0(CLBLL_R_X71Y118_SLICE_X107Y118_BO6),
.I1(CLBLL_R_X71Y118_SLICE_X107Y118_AO6),
.O(CLBLL_R_X71Y118_SLICE_X107Y118_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y118_SLICE_X107Y118_MUXF7B (
.I0(CLBLL_R_X71Y118_SLICE_X107Y118_DO6),
.I1(CLBLL_R_X71Y118_SLICE_X107Y118_CO6),
.O(CLBLL_R_X71Y118_SLICE_X107Y118_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X71Y118_SLICE_X107Y118_MUXF8 (
.I0(CLBLL_R_X71Y118_SLICE_X107Y118_F7BMUX_O),
.I1(CLBLL_R_X71Y118_SLICE_X107Y118_F7AMUX_O),
.O(CLBLL_R_X71Y118_SLICE_X107Y118_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLL_R_X71Y119_SLICE_X106Y119_AO6),
.Q(CLBLL_R_X71Y119_SLICE_X106Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h689e59a195636e96)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_DLUT (
.I0(CLBLM_L_X74Y117_SLICE_X113Y117_DO6),
.I1(CLBLL_R_X75Y120_SLICE_X115Y120_CO6),
.I2(CLBLL_R_X73Y116_SLICE_X110Y116_CO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_CO6),
.I4(CLBLM_L_X72Y116_SLICE_X108Y116_DO6),
.I5(CLBLM_L_X74Y117_SLICE_X113Y117_CO6),
.O5(CLBLL_R_X71Y119_SLICE_X106Y119_DO5),
.O6(CLBLL_R_X71Y119_SLICE_X106Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he41b38c61ed53c2b)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_CLUT (
.I0(CLBLM_L_X74Y117_SLICE_X113Y117_DO6),
.I1(CLBLL_R_X75Y120_SLICE_X115Y120_CO6),
.I2(CLBLL_R_X73Y116_SLICE_X110Y116_CO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_CO6),
.I4(CLBLM_L_X72Y116_SLICE_X108Y116_DO6),
.I5(CLBLM_L_X74Y117_SLICE_X113Y117_CO6),
.O5(CLBLL_R_X71Y119_SLICE_X106Y119_CO5),
.O6(CLBLL_R_X71Y119_SLICE_X106Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4c34d781bacd662)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_BLUT (
.I0(CLBLM_L_X72Y116_SLICE_X108Y116_DO6),
.I1(CLBLM_L_X74Y117_SLICE_X113Y117_CO6),
.I2(CLBLL_R_X73Y116_SLICE_X110Y116_CO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_CO6),
.I4(CLBLM_L_X74Y117_SLICE_X113Y117_DO6),
.I5(CLBLL_R_X75Y120_SLICE_X115Y120_CO6),
.O5(CLBLL_R_X71Y119_SLICE_X106Y119_BO5),
.O6(CLBLL_R_X71Y119_SLICE_X106Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ccf5cca0)
  ) CLBLL_R_X71Y119_SLICE_X106Y119_ALUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I1(RIOB33_X105Y151_IOB_X1Y151_I),
.I2(CLBLL_R_X71Y119_SLICE_X106Y119_AQ),
.I3(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I4(CLBLM_L_X70Y119_SLICE_X104Y119_AQ),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.O5(CLBLL_R_X71Y119_SLICE_X106Y119_AO5),
.O6(CLBLL_R_X71Y119_SLICE_X106Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fcacaf000caca)
  ) CLBLL_R_X71Y119_SLICE_X107Y119_DLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.O5(CLBLL_R_X71Y119_SLICE_X107Y119_DO5),
.O6(CLBLL_R_X71Y119_SLICE_X107Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefece3e02f2c2320)
  ) CLBLL_R_X71Y119_SLICE_X107Y119_CLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I5(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.O5(CLBLL_R_X71Y119_SLICE_X107Y119_CO5),
.O6(CLBLL_R_X71Y119_SLICE_X107Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cfcfc0c0)
  ) CLBLL_R_X71Y119_SLICE_X107Y119_BLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X71Y119_SLICE_X107Y119_BO5),
.O6(CLBLL_R_X71Y119_SLICE_X107Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff00cccc)
  ) CLBLL_R_X71Y119_SLICE_X107Y119_ALUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I3(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X71Y119_SLICE_X107Y119_AO5),
.O6(CLBLL_R_X71Y119_SLICE_X107Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y119_SLICE_X107Y119_MUXF7A (
.I0(CLBLL_R_X71Y119_SLICE_X107Y119_BO6),
.I1(CLBLL_R_X71Y119_SLICE_X107Y119_AO6),
.O(CLBLL_R_X71Y119_SLICE_X107Y119_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y119_SLICE_X107Y119_MUXF7B (
.I0(CLBLL_R_X71Y119_SLICE_X107Y119_DO6),
.I1(CLBLL_R_X71Y119_SLICE_X107Y119_CO6),
.O(CLBLL_R_X71Y119_SLICE_X107Y119_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf85d58ada80d08)
  ) CLBLL_R_X71Y120_SLICE_X106Y120_DLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I4(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.O5(CLBLL_R_X71Y120_SLICE_X106Y120_DO5),
.O6(CLBLL_R_X71Y120_SLICE_X106Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ff55aa00)
  ) CLBLL_R_X71Y120_SLICE_X106Y120_CLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X71Y120_SLICE_X106Y120_CO5),
.O6(CLBLL_R_X71Y120_SLICE_X106Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccff00f0f0)
  ) CLBLL_R_X71Y120_SLICE_X106Y120_BLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I1(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X71Y120_SLICE_X106Y120_BO5),
.O6(CLBLL_R_X71Y120_SLICE_X106Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaccccf0f0)
  ) CLBLL_R_X71Y120_SLICE_X106Y120_ALUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X71Y120_SLICE_X106Y120_AO5),
.O6(CLBLL_R_X71Y120_SLICE_X106Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y120_SLICE_X106Y120_MUXF7A (
.I0(CLBLL_R_X71Y120_SLICE_X106Y120_BO6),
.I1(CLBLL_R_X71Y120_SLICE_X106Y120_AO6),
.O(CLBLL_R_X71Y120_SLICE_X106Y120_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y120_SLICE_X106Y120_MUXF7B (
.I0(CLBLL_R_X71Y120_SLICE_X106Y120_DO6),
.I1(CLBLL_R_X71Y120_SLICE_X106Y120_CO6),
.O(CLBLL_R_X71Y120_SLICE_X106Y120_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96a5c53259c669ad)
  ) CLBLL_R_X71Y120_SLICE_X107Y120_DLUT (
.I0(CLBLL_R_X71Y120_SLICE_X107Y120_AO6),
.I1(CLBLL_R_X71Y122_SLICE_X106Y122_AO6),
.I2(CLBLL_R_X73Y120_SLICE_X111Y120_DO6),
.I3(CLBLM_L_X72Y120_SLICE_X108Y120_DO6),
.I4(CLBLL_R_X73Y120_SLICE_X111Y120_CO6),
.I5(CLBLM_L_X74Y120_SLICE_X113Y120_AO6),
.O5(CLBLL_R_X71Y120_SLICE_X107Y120_DO5),
.O6(CLBLL_R_X71Y120_SLICE_X107Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd263691bd4e42b)
  ) CLBLL_R_X71Y120_SLICE_X107Y120_CLUT (
.I0(CLBLL_R_X71Y120_SLICE_X107Y120_AO6),
.I1(CLBLM_L_X74Y120_SLICE_X113Y120_AO6),
.I2(CLBLM_L_X72Y120_SLICE_X108Y120_DO6),
.I3(CLBLL_R_X71Y122_SLICE_X106Y122_AO6),
.I4(CLBLL_R_X73Y120_SLICE_X111Y120_CO6),
.I5(CLBLL_R_X73Y120_SLICE_X111Y120_DO6),
.O5(CLBLL_R_X71Y120_SLICE_X107Y120_CO5),
.O6(CLBLL_R_X71Y120_SLICE_X107Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5c31af0788f671c)
  ) CLBLL_R_X71Y120_SLICE_X107Y120_BLUT (
.I0(CLBLL_R_X73Y120_SLICE_X111Y120_CO6),
.I1(CLBLM_L_X74Y120_SLICE_X113Y120_AO6),
.I2(CLBLM_L_X72Y120_SLICE_X108Y120_DO6),
.I3(CLBLL_R_X73Y120_SLICE_X111Y120_DO6),
.I4(CLBLL_R_X71Y120_SLICE_X107Y120_AO6),
.I5(CLBLL_R_X71Y122_SLICE_X106Y122_AO6),
.O5(CLBLL_R_X71Y120_SLICE_X107Y120_BO5),
.O6(CLBLL_R_X71Y120_SLICE_X107Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h569a5555569aaaaa)
  ) CLBLL_R_X71Y120_SLICE_X107Y120_ALUT (
.I0(CLBLM_L_X70Y127_SLICE_X104Y127_DO6),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLL_R_X71Y119_SLICE_X107Y119_F7BMUX_O),
.I3(CLBLL_R_X71Y120_SLICE_X106Y120_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLM_L_X72Y120_SLICE_X109Y120_F8MUX_O),
.O5(CLBLL_R_X71Y120_SLICE_X107Y120_AO5),
.O6(CLBLL_R_X71Y120_SLICE_X107Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcee223030ee22)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_DLUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I1(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.O5(CLBLL_R_X71Y121_SLICE_X106Y121_DO5),
.O6(CLBLL_R_X71Y121_SLICE_X106Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf83b38cbc80b08)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_CLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I1(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.O5(CLBLL_R_X71Y121_SLICE_X106Y121_CO5),
.O6(CLBLL_R_X71Y121_SLICE_X106Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaffca0fcaf0ca00)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_BLUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.O5(CLBLL_R_X71Y121_SLICE_X106Y121_BO5),
.O6(CLBLL_R_X71Y121_SLICE_X106Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeef5a04444f5a0)
  ) CLBLL_R_X71Y121_SLICE_X106Y121_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.O5(CLBLL_R_X71Y121_SLICE_X106Y121_AO5),
.O6(CLBLL_R_X71Y121_SLICE_X106Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y121_SLICE_X106Y121_MUXF7A (
.I0(CLBLL_R_X71Y121_SLICE_X106Y121_BO6),
.I1(CLBLL_R_X71Y121_SLICE_X106Y121_AO6),
.O(CLBLL_R_X71Y121_SLICE_X106Y121_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y121_SLICE_X106Y121_MUXF7B (
.I0(CLBLL_R_X71Y121_SLICE_X106Y121_DO6),
.I1(CLBLL_R_X71Y121_SLICE_X106Y121_CO6),
.O(CLBLL_R_X71Y121_SLICE_X106Y121_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cafaffc0ca0a0)
  ) CLBLL_R_X71Y121_SLICE_X107Y121_DLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.O5(CLBLL_R_X71Y121_SLICE_X107Y121_DO5),
.O6(CLBLL_R_X71Y121_SLICE_X107Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cfcfafa0c0c0)
  ) CLBLL_R_X71Y121_SLICE_X107Y121_CLUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.O5(CLBLL_R_X71Y121_SLICE_X107Y121_CO5),
.O6(CLBLL_R_X71Y121_SLICE_X107Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaef4a45e0e5404)
  ) CLBLL_R_X71Y121_SLICE_X107Y121_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I4(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.O5(CLBLL_R_X71Y121_SLICE_X107Y121_BO5),
.O6(CLBLL_R_X71Y121_SLICE_X107Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaf0f0ff00)
  ) CLBLL_R_X71Y121_SLICE_X107Y121_ALUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLL_R_X71Y121_SLICE_X107Y121_AO5),
.O6(CLBLL_R_X71Y121_SLICE_X107Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y121_SLICE_X107Y121_MUXF7A (
.I0(CLBLL_R_X71Y121_SLICE_X107Y121_BO6),
.I1(CLBLL_R_X71Y121_SLICE_X107Y121_AO6),
.O(CLBLL_R_X71Y121_SLICE_X107Y121_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y121_SLICE_X107Y121_MUXF7B (
.I0(CLBLL_R_X71Y121_SLICE_X107Y121_DO6),
.I1(CLBLL_R_X71Y121_SLICE_X107Y121_CO6),
.O(CLBLL_R_X71Y121_SLICE_X107Y121_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X71Y121_SLICE_X107Y121_MUXF8 (
.I0(CLBLL_R_X71Y121_SLICE_X107Y121_F7BMUX_O),
.I1(CLBLL_R_X71Y121_SLICE_X107Y121_F7AMUX_O),
.O(CLBLL_R_X71Y121_SLICE_X107Y121_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y122_SLICE_X106Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y122_SLICE_X106Y122_DO5),
.O6(CLBLL_R_X71Y122_SLICE_X106Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y122_SLICE_X106Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y122_SLICE_X106Y122_CO5),
.O6(CLBLL_R_X71Y122_SLICE_X106Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y122_SLICE_X106Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y122_SLICE_X106Y122_BO5),
.O6(CLBLL_R_X71Y122_SLICE_X106Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05faf50a35ca35ca)
  ) CLBLL_R_X71Y122_SLICE_X106Y122_ALUT (
.I0(CLBLL_R_X71Y121_SLICE_X107Y121_F8MUX_O),
.I1(CLBLL_R_X71Y121_SLICE_X106Y121_F7AMUX_O),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(CLBLL_L_X2Y124_SLICE_X0Y124_CO6),
.I4(CLBLL_R_X71Y121_SLICE_X106Y121_F7BMUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X71Y122_SLICE_X106Y122_AO5),
.O6(CLBLL_R_X71Y122_SLICE_X106Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y122_SLICE_X107Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y122_SLICE_X107Y122_DO5),
.O6(CLBLL_R_X71Y122_SLICE_X107Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y122_SLICE_X107Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y122_SLICE_X107Y122_CO5),
.O6(CLBLL_R_X71Y122_SLICE_X107Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y122_SLICE_X107Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y122_SLICE_X107Y122_BO5),
.O6(CLBLL_R_X71Y122_SLICE_X107Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y122_SLICE_X107Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y122_SLICE_X107Y122_AO5),
.O6(CLBLL_R_X71Y122_SLICE_X107Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9679626c79868697)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_DLUT (
.I0(CLBLL_R_X71Y127_SLICE_X107Y127_AO6),
.I1(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I2(CLBLL_R_X71Y125_SLICE_X107Y125_DO6),
.I3(CLBLM_L_X72Y128_SLICE_X108Y128_CO6),
.I4(CLBLL_R_X71Y126_SLICE_X107Y126_DO6),
.I5(CLBLL_R_X75Y125_SLICE_X115Y125_DO6),
.O5(CLBLL_R_X71Y125_SLICE_X106Y125_DO5),
.O6(CLBLL_R_X71Y125_SLICE_X106Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha96d96165ae4659a)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_CLUT (
.I0(CLBLL_R_X71Y127_SLICE_X107Y127_AO6),
.I1(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I2(CLBLL_R_X71Y125_SLICE_X107Y125_DO6),
.I3(CLBLM_L_X72Y128_SLICE_X108Y128_CO6),
.I4(CLBLL_R_X71Y126_SLICE_X107Y126_DO6),
.I5(CLBLL_R_X75Y125_SLICE_X115Y125_DO6),
.O5(CLBLL_R_X71Y125_SLICE_X106Y125_CO5),
.O6(CLBLL_R_X71Y125_SLICE_X106Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h64bf39c78ba0d429)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_BLUT (
.I0(CLBLL_R_X71Y126_SLICE_X107Y126_DO6),
.I1(CLBLL_R_X71Y125_SLICE_X107Y125_DO6),
.I2(CLBLL_R_X71Y127_SLICE_X107Y127_AO6),
.I3(CLBLL_R_X75Y125_SLICE_X115Y125_DO6),
.I4(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I5(CLBLM_L_X72Y128_SLICE_X108Y128_CO6),
.O5(CLBLL_R_X71Y125_SLICE_X106Y125_BO5),
.O6(CLBLL_R_X71Y125_SLICE_X106Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6919d9a69649a676)
  ) CLBLL_R_X71Y125_SLICE_X106Y125_ALUT (
.I0(CLBLL_R_X71Y126_SLICE_X107Y126_DO6),
.I1(CLBLL_R_X71Y125_SLICE_X107Y125_DO6),
.I2(CLBLL_R_X71Y127_SLICE_X107Y127_AO6),
.I3(CLBLL_R_X75Y125_SLICE_X115Y125_DO6),
.I4(CLBLL_R_X71Y125_SLICE_X107Y125_CO6),
.I5(CLBLM_L_X72Y128_SLICE_X108Y128_CO6),
.O5(CLBLL_R_X71Y125_SLICE_X106Y125_AO5),
.O6(CLBLL_R_X71Y125_SLICE_X106Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h101fd0dfefe02f20)
  ) CLBLL_R_X71Y125_SLICE_X107Y125_DLUT (
.I0(CLBLM_L_X72Y125_SLICE_X108Y125_F7BMUX_O),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(CLBLM_L_X72Y125_SLICE_X109Y125_F8MUX_O),
.I4(CLBLM_L_X72Y124_SLICE_X108Y124_F7AMUX_O),
.I5(CLBLM_L_X70Y128_SLICE_X104Y128_BO6),
.O5(CLBLL_R_X71Y125_SLICE_X107Y125_DO5),
.O6(CLBLL_R_X71Y125_SLICE_X107Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h556699aa5a5a5a5a)
  ) CLBLL_R_X71Y125_SLICE_X107Y125_CLUT (
.I0(CLBLM_L_X56Y116_SLICE_X84Y116_CO6),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLL_R_X73Y125_SLICE_X110Y125_F8MUX_O),
.I3(CLBLL_R_X71Y125_SLICE_X107Y125_F7AMUX_O),
.I4(CLBLM_L_X72Y125_SLICE_X108Y125_F7AMUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLL_R_X71Y125_SLICE_X107Y125_CO5),
.O6(CLBLL_R_X71Y125_SLICE_X107Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbf3bbc088f388c0)
  ) CLBLL_R_X71Y125_SLICE_X107Y125_BLUT (
.I0(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.O5(CLBLL_R_X71Y125_SLICE_X107Y125_BO5),
.O6(CLBLL_R_X71Y125_SLICE_X107Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3eef322c0eec022)
  ) CLBLL_R_X71Y125_SLICE_X107Y125_ALUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I5(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.O5(CLBLL_R_X71Y125_SLICE_X107Y125_AO5),
.O6(CLBLL_R_X71Y125_SLICE_X107Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y125_SLICE_X107Y125_MUXF7A (
.I0(CLBLL_R_X71Y125_SLICE_X107Y125_BO6),
.I1(CLBLL_R_X71Y125_SLICE_X107Y125_AO6),
.O(CLBLL_R_X71Y125_SLICE_X107Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y126_SLICE_X106Y126_DO5),
.O6(CLBLL_R_X71Y126_SLICE_X106Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y126_SLICE_X106Y126_CO5),
.O6(CLBLL_R_X71Y126_SLICE_X106Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h652ee992295592eb)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_BLUT (
.I0(CLBLL_R_X75Y125_SLICE_X115Y125_CO6),
.I1(CLBLL_R_X75Y125_SLICE_X114Y125_CO6),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_CO6),
.I3(CLBLM_L_X72Y124_SLICE_X108Y124_CO6),
.I4(CLBLM_L_X74Y125_SLICE_X112Y125_CO6),
.I5(CLBLL_R_X73Y127_SLICE_X111Y127_CO6),
.O5(CLBLL_R_X71Y126_SLICE_X106Y126_BO5),
.O6(CLBLL_R_X71Y126_SLICE_X106Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd6792a9543aeb642)
  ) CLBLL_R_X71Y126_SLICE_X106Y126_ALUT (
.I0(CLBLL_R_X75Y125_SLICE_X115Y125_CO6),
.I1(CLBLL_R_X75Y125_SLICE_X114Y125_CO6),
.I2(CLBLL_R_X71Y126_SLICE_X107Y126_CO6),
.I3(CLBLL_R_X73Y127_SLICE_X111Y127_CO6),
.I4(CLBLM_L_X74Y125_SLICE_X112Y125_CO6),
.I5(CLBLM_L_X72Y124_SLICE_X108Y124_CO6),
.O5(CLBLL_R_X71Y126_SLICE_X106Y126_AO5),
.O6(CLBLL_R_X71Y126_SLICE_X106Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa66665a5a6666)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_DLUT (
.I0(CLBLL_R_X71Y128_SLICE_X106Y128_CO6),
.I1(CLBLM_L_X72Y126_SLICE_X108Y126_F8MUX_O),
.I2(CLBLM_L_X72Y126_SLICE_X109Y126_F7BMUX_O),
.I3(CLBLL_R_X71Y126_SLICE_X107Y126_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X71Y126_SLICE_X107Y126_DO5),
.O6(CLBLL_R_X71Y126_SLICE_X107Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55330f0faaccf0f0)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_CLUT (
.I0(CLBLL_R_X73Y126_SLICE_X111Y126_F7BMUX_O),
.I1(CLBLM_L_X72Y126_SLICE_X109Y126_F7AMUX_O),
.I2(CLBLL_R_X73Y126_SLICE_X110Y126_F8MUX_O),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.O5(CLBLL_R_X71Y126_SLICE_X107Y126_CO5),
.O6(CLBLL_R_X71Y126_SLICE_X107Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2ff33e2e2cc00)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_BLUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.O5(CLBLL_R_X71Y126_SLICE_X107Y126_BO5),
.O6(CLBLL_R_X71Y126_SLICE_X107Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0aaffccf0aa00)
  ) CLBLL_R_X71Y126_SLICE_X107Y126_ALUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I2(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.O5(CLBLL_R_X71Y126_SLICE_X107Y126_AO5),
.O6(CLBLL_R_X71Y126_SLICE_X107Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X71Y126_SLICE_X107Y126_MUXF7A (
.I0(CLBLL_R_X71Y126_SLICE_X107Y126_BO6),
.I1(CLBLL_R_X71Y126_SLICE_X107Y126_AO6),
.O(CLBLL_R_X71Y126_SLICE_X107Y126_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y127_SLICE_X106Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X106Y127_DO5),
.O6(CLBLL_R_X71Y127_SLICE_X106Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y127_SLICE_X106Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X106Y127_CO5),
.O6(CLBLL_R_X71Y127_SLICE_X106Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hce23355a37d80a6d)
  ) CLBLL_R_X71Y127_SLICE_X106Y127_BLUT (
.I0(CLBLL_R_X73Y127_SLICE_X111Y127_CO6),
.I1(CLBLM_L_X72Y124_SLICE_X108Y124_CO6),
.I2(CLBLM_L_X74Y125_SLICE_X112Y125_CO6),
.I3(CLBLL_R_X75Y125_SLICE_X115Y125_CO6),
.I4(CLBLL_R_X75Y125_SLICE_X114Y125_CO6),
.I5(CLBLL_R_X71Y126_SLICE_X107Y126_CO6),
.O5(CLBLL_R_X71Y127_SLICE_X106Y127_BO5),
.O6(CLBLL_R_X71Y127_SLICE_X106Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h998786764e31962f)
  ) CLBLL_R_X71Y127_SLICE_X106Y127_ALUT (
.I0(CLBLL_R_X73Y127_SLICE_X111Y127_CO6),
.I1(CLBLM_L_X72Y124_SLICE_X108Y124_CO6),
.I2(CLBLM_L_X74Y125_SLICE_X112Y125_CO6),
.I3(CLBLL_R_X75Y125_SLICE_X115Y125_CO6),
.I4(CLBLL_R_X75Y125_SLICE_X114Y125_CO6),
.I5(CLBLL_R_X71Y126_SLICE_X107Y126_CO6),
.O5(CLBLL_R_X71Y127_SLICE_X106Y127_AO5),
.O6(CLBLL_R_X71Y127_SLICE_X106Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X107Y127_DO5),
.O6(CLBLL_R_X71Y127_SLICE_X107Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X107Y127_CO5),
.O6(CLBLL_R_X71Y127_SLICE_X107Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y127_SLICE_X107Y127_BO5),
.O6(CLBLL_R_X71Y127_SLICE_X107Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05f53535fa0acaca)
  ) CLBLL_R_X71Y127_SLICE_X107Y127_ALUT (
.I0(CLBLM_L_X72Y127_SLICE_X109Y127_F8MUX_O),
.I1(CLBLM_L_X72Y127_SLICE_X108Y127_F7AMUX_O),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(CLBLM_L_X72Y127_SLICE_X108Y127_F7BMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_L_X2Y118_SLICE_X0Y118_CO6),
.O5(CLBLL_R_X71Y127_SLICE_X107Y127_AO5),
.O6(CLBLL_R_X71Y127_SLICE_X107Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLL_R_X71Y128_SLICE_X106Y128_CO6),
.Q(CLBLL_R_X71Y128_SLICE_X106Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLL_R_X71Y128_SLICE_X106Y128_AO6),
.Q(CLBLL_R_X71Y128_SLICE_X106Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X106Y128_DO5),
.O6(CLBLL_R_X71Y128_SLICE_X106Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f1f1e0e0)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_CLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I2(CLBLL_R_X71Y128_SLICE_X106Y128_AQ),
.I3(RIOB33_X105Y155_IOB_X1Y155_I),
.I4(CLBLL_R_X71Y128_SLICE_X106Y128_BQ),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLL_R_X71Y128_SLICE_X106Y128_CO5),
.O6(CLBLL_R_X71Y128_SLICE_X106Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0ccf0ccf0aa)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_BLUT (
.I0(RIOB33_X105Y153_IOB_X1Y154_I),
.I1(CLBLL_R_X71Y128_SLICE_X106Y128_BQ),
.I2(CLBLL_R_X71Y128_SLICE_X106Y128_AQ),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X71Y128_SLICE_X106Y128_BO5),
.O6(CLBLL_R_X71Y128_SLICE_X106Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00e1ff1e0)
  ) CLBLL_R_X71Y128_SLICE_X106Y128_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLL_R_X71Y128_SLICE_X106Y128_AQ),
.I3(CLBLL_R_X71Y128_SLICE_X106Y128_BO6),
.I4(CLBLL_R_X71Y127_SLICE_X106Y127_BO6),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLL_R_X71Y128_SLICE_X106Y128_AO5),
.O6(CLBLL_R_X71Y128_SLICE_X106Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X107Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X107Y128_DO5),
.O6(CLBLL_R_X71Y128_SLICE_X107Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X107Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X107Y128_CO5),
.O6(CLBLL_R_X71Y128_SLICE_X107Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X107Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X107Y128_BO5),
.O6(CLBLL_R_X71Y128_SLICE_X107Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y128_SLICE_X107Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y128_SLICE_X107Y128_AO5),
.O6(CLBLL_R_X71Y128_SLICE_X107Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X106Y129_DO5),
.O6(CLBLL_R_X71Y129_SLICE_X106Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X106Y129_CO5),
.O6(CLBLL_R_X71Y129_SLICE_X106Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X106Y129_BO5),
.O6(CLBLL_R_X71Y129_SLICE_X106Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf26989a72c26799c)
  ) CLBLL_R_X71Y129_SLICE_X106Y129_ALUT (
.I0(CLBLL_R_X73Y129_SLICE_X110Y129_CO6),
.I1(CLBLL_R_X75Y127_SLICE_X114Y127_CO6),
.I2(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I3(CLBLM_L_X74Y128_SLICE_X112Y128_CO6),
.I4(CLBLM_L_X72Y128_SLICE_X109Y128_DO6),
.I5(CLBLM_L_X72Y128_SLICE_X109Y128_CO6),
.O5(CLBLL_R_X71Y129_SLICE_X106Y129_AO5),
.O6(CLBLL_R_X71Y129_SLICE_X106Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X107Y129_DO5),
.O6(CLBLL_R_X71Y129_SLICE_X107Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X107Y129_CO5),
.O6(CLBLL_R_X71Y129_SLICE_X107Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X107Y129_BO5),
.O6(CLBLL_R_X71Y129_SLICE_X107Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X71Y129_SLICE_X107Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X71Y129_SLICE_X107Y129_AO5),
.O6(CLBLL_R_X71Y129_SLICE_X107Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLL_R_X71Y131_SLICE_X106Y131_CO6),
.Q(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLL_R_X71Y131_SLICE_X106Y131_AO6),
.Q(CLBLL_R_X71Y131_SLICE_X106Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hac1a63c595c7d869)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_DLUT (
.I0(CLBLM_L_X72Y128_SLICE_X109Y128_DO6),
.I1(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I2(CLBLL_R_X73Y129_SLICE_X110Y129_CO6),
.I3(CLBLM_L_X74Y128_SLICE_X112Y128_CO6),
.I4(CLBLL_R_X75Y127_SLICE_X114Y127_CO6),
.I5(CLBLM_L_X72Y128_SLICE_X109Y128_CO6),
.O5(CLBLL_R_X71Y131_SLICE_X106Y131_DO5),
.O6(CLBLL_R_X71Y131_SLICE_X106Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfdfcec30313020)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_CLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I1(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I2(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I4(CLBLL_R_X71Y131_SLICE_X106Y131_BQ),
.I5(RIOB33_X105Y163_IOB_X1Y163_I),
.O5(CLBLL_R_X71Y131_SLICE_X106Y131_CO5),
.O6(CLBLL_R_X71Y131_SLICE_X106Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e2e2e2e2f3c0)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_BLUT (
.I0(CLBLL_R_X71Y131_SLICE_X106Y131_BQ),
.I1(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I2(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I3(RIOB33_X105Y161_IOB_X1Y162_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X71Y131_SLICE_X106Y131_BO5),
.O6(CLBLL_R_X71Y131_SLICE_X106Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a596a)
  ) CLBLL_R_X71Y131_SLICE_X106Y131_ALUT (
.I0(CLBLL_R_X71Y131_SLICE_X106Y131_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(CLBLL_R_X71Y131_SLICE_X106Y131_AQ),
.I3(CLBLL_R_X71Y131_SLICE_X106Y131_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X71Y131_SLICE_X106Y131_AO5),
.O6(CLBLL_R_X71Y131_SLICE_X106Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLL_R_X71Y131_SLICE_X107Y131_DO6),
.Q(CLBLL_R_X71Y131_SLICE_X107Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLL_R_X71Y131_SLICE_X107Y131_BO6),
.Q(CLBLL_R_X71Y131_SLICE_X107Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X72Y131_SLICE_X108Y131_AO6),
.Q(CLBLL_R_X71Y131_SLICE_X107Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffee1100)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_DLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I2(RIOB33_X105Y157_IOB_X1Y157_I),
.I3(CLBLL_R_X71Y131_SLICE_X107Y131_BQ),
.I4(CLBLL_R_X71Y131_SLICE_X107Y131_AQ),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLL_R_X71Y131_SLICE_X107Y131_DO5),
.O6(CLBLL_R_X71Y131_SLICE_X107Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fe987610)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_CLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(RIOB33_X105Y155_IOB_X1Y156_I),
.I3(CLBLL_R_X71Y131_SLICE_X107Y131_BQ),
.I4(CLBLL_R_X71Y131_SLICE_X107Y131_AQ),
.I5(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.O5(CLBLL_R_X71Y131_SLICE_X107Y131_CO5),
.O6(CLBLL_R_X71Y131_SLICE_X107Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h666666666663666c)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_BLUT (
.I0(CLBLL_R_X71Y131_SLICE_X107Y131_AQ),
.I1(CLBLM_L_X72Y131_SLICE_X108Y131_CO6),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(LIOB33_X0Y79_IOB_X0Y80_I),
.I4(CLBLL_R_X71Y131_SLICE_X107Y131_CO6),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X71Y131_SLICE_X107Y131_BO5),
.O6(CLBLL_R_X71Y131_SLICE_X107Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aafcaa30)
  ) CLBLL_R_X71Y131_SLICE_X107Y131_ALUT (
.I0(RIOB33_X105Y171_IOB_X1Y171_I),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I2(CLBLL_R_X71Y131_SLICE_X107Y131_CQ),
.I3(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I4(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.O5(CLBLL_R_X71Y131_SLICE_X107Y131_AO5),
.O6(CLBLL_R_X71Y131_SLICE_X107Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaffca0fcaf0ca00)
  ) CLBLL_R_X73Y114_SLICE_X110Y114_DLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.O5(CLBLL_R_X73Y114_SLICE_X110Y114_DO5),
.O6(CLBLL_R_X73Y114_SLICE_X110Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcaf0caffca00ca0)
  ) CLBLL_R_X73Y114_SLICE_X110Y114_CLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I1(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.O5(CLBLL_R_X73Y114_SLICE_X110Y114_CO5),
.O6(CLBLL_R_X73Y114_SLICE_X110Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef4fea4ae545e040)
  ) CLBLL_R_X73Y114_SLICE_X110Y114_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.O5(CLBLL_R_X73Y114_SLICE_X110Y114_BO5),
.O6(CLBLL_R_X73Y114_SLICE_X110Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacafff00f00)
  ) CLBLL_R_X73Y114_SLICE_X110Y114_ALUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I4(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y114_SLICE_X110Y114_AO5),
.O6(CLBLL_R_X73Y114_SLICE_X110Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y114_SLICE_X110Y114_MUXF7A (
.I0(CLBLL_R_X73Y114_SLICE_X110Y114_BO6),
.I1(CLBLL_R_X73Y114_SLICE_X110Y114_AO6),
.O(CLBLL_R_X73Y114_SLICE_X110Y114_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y114_SLICE_X110Y114_MUXF7B (
.I0(CLBLL_R_X73Y114_SLICE_X110Y114_DO6),
.I1(CLBLL_R_X73Y114_SLICE_X110Y114_CO6),
.O(CLBLL_R_X73Y114_SLICE_X110Y114_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y114_SLICE_X110Y114_MUXF8 (
.I0(CLBLL_R_X73Y114_SLICE_X110Y114_F7BMUX_O),
.I1(CLBLL_R_X73Y114_SLICE_X110Y114_F7AMUX_O),
.O(CLBLL_R_X73Y114_SLICE_X110Y114_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y114_SLICE_X111Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y114_SLICE_X111Y114_DO5),
.O6(CLBLL_R_X73Y114_SLICE_X111Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y114_SLICE_X111Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y114_SLICE_X111Y114_CO5),
.O6(CLBLL_R_X73Y114_SLICE_X111Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y114_SLICE_X111Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y114_SLICE_X111Y114_BO5),
.O6(CLBLL_R_X73Y114_SLICE_X111Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y114_SLICE_X111Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y114_SLICE_X111Y114_AO5),
.O6(CLBLL_R_X73Y114_SLICE_X111Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y115_SLICE_X110Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y115_SLICE_X110Y115_DO5),
.O6(CLBLL_R_X73Y115_SLICE_X110Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05278daffad87250)
  ) CLBLL_R_X73Y115_SLICE_X110Y115_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLL_R_X73Y115_SLICE_X111Y115_F8MUX_O),
.I3(CLBLL_R_X73Y115_SLICE_X110Y115_F7AMUX_O),
.I4(CLBLM_L_X72Y115_SLICE_X109Y115_F7AMUX_O),
.I5(CLBLL_R_X71Y119_SLICE_X106Y119_AO6),
.O5(CLBLL_R_X73Y115_SLICE_X110Y115_CO5),
.O6(CLBLL_R_X73Y115_SLICE_X110Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddf5dda088f588a0)
  ) CLBLL_R_X73Y115_SLICE_X110Y115_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.O5(CLBLL_R_X73Y115_SLICE_X110Y115_BO5),
.O6(CLBLL_R_X73Y115_SLICE_X110Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4ffe455e4aae400)
  ) CLBLL_R_X73Y115_SLICE_X110Y115_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I5(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.O5(CLBLL_R_X73Y115_SLICE_X110Y115_AO5),
.O6(CLBLL_R_X73Y115_SLICE_X110Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y115_SLICE_X110Y115_MUXF7A (
.I0(CLBLL_R_X73Y115_SLICE_X110Y115_BO6),
.I1(CLBLL_R_X73Y115_SLICE_X110Y115_AO6),
.O(CLBLL_R_X73Y115_SLICE_X110Y115_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcee30eefc223022)
  ) CLBLL_R_X73Y115_SLICE_X111Y115_DLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.O5(CLBLL_R_X73Y115_SLICE_X111Y115_DO5),
.O6(CLBLL_R_X73Y115_SLICE_X111Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaccf0ccf0)
  ) CLBLL_R_X73Y115_SLICE_X111Y115_CLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y115_SLICE_X111Y115_CO5),
.O6(CLBLL_R_X73Y115_SLICE_X111Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ff55aa00)
  ) CLBLL_R_X73Y115_SLICE_X111Y115_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I3(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X73Y115_SLICE_X111Y115_BO5),
.O6(CLBLL_R_X73Y115_SLICE_X111Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0eeeef5a04444)
  ) CLBLL_R_X73Y115_SLICE_X111Y115_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.O5(CLBLL_R_X73Y115_SLICE_X111Y115_AO5),
.O6(CLBLL_R_X73Y115_SLICE_X111Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y115_SLICE_X111Y115_MUXF7A (
.I0(CLBLL_R_X73Y115_SLICE_X111Y115_BO6),
.I1(CLBLL_R_X73Y115_SLICE_X111Y115_AO6),
.O(CLBLL_R_X73Y115_SLICE_X111Y115_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y115_SLICE_X111Y115_MUXF7B (
.I0(CLBLL_R_X73Y115_SLICE_X111Y115_DO6),
.I1(CLBLL_R_X73Y115_SLICE_X111Y115_CO6),
.O(CLBLL_R_X73Y115_SLICE_X111Y115_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y115_SLICE_X111Y115_MUXF8 (
.I0(CLBLL_R_X73Y115_SLICE_X111Y115_F7BMUX_O),
.I1(CLBLL_R_X73Y115_SLICE_X111Y115_F7AMUX_O),
.O(CLBLL_R_X73Y115_SLICE_X111Y115_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y116_SLICE_X110Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y116_SLICE_X110Y116_DO5),
.O6(CLBLL_R_X73Y116_SLICE_X110Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h569a569a56569a9a)
  ) CLBLL_R_X73Y116_SLICE_X110Y116_CLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(CLBLL_R_X73Y116_SLICE_X111Y116_F8MUX_O),
.I3(CLBLL_R_X73Y116_SLICE_X110Y116_F7AMUX_O),
.I4(CLBLM_L_X72Y116_SLICE_X109Y116_F7BMUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X73Y116_SLICE_X110Y116_CO5),
.O6(CLBLL_R_X73Y116_SLICE_X110Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fcfc0c0c)
  ) CLBLL_R_X73Y116_SLICE_X110Y116_BLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y116_SLICE_X110Y116_BO5),
.O6(CLBLL_R_X73Y116_SLICE_X110Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd855d8aad800d8)
  ) CLBLL_R_X73Y116_SLICE_X110Y116_ALUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.O5(CLBLL_R_X73Y116_SLICE_X110Y116_AO5),
.O6(CLBLL_R_X73Y116_SLICE_X110Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y116_SLICE_X110Y116_MUXF7A (
.I0(CLBLL_R_X73Y116_SLICE_X110Y116_BO6),
.I1(CLBLL_R_X73Y116_SLICE_X110Y116_AO6),
.O(CLBLL_R_X73Y116_SLICE_X110Y116_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfafafc0c0a0a)
  ) CLBLL_R_X73Y116_SLICE_X111Y116_DLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.O5(CLBLL_R_X73Y116_SLICE_X111Y116_DO5),
.O6(CLBLL_R_X73Y116_SLICE_X111Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccb8b83300b8b8)
  ) CLBLL_R_X73Y116_SLICE_X111Y116_CLUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.O5(CLBLL_R_X73Y116_SLICE_X111Y116_CO5),
.O6(CLBLL_R_X73Y116_SLICE_X111Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcee30eefc223022)
  ) CLBLL_R_X73Y116_SLICE_X111Y116_BLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.O5(CLBLL_R_X73Y116_SLICE_X111Y116_BO5),
.O6(CLBLL_R_X73Y116_SLICE_X111Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbcbf8c83b0b3808)
  ) CLBLL_R_X73Y116_SLICE_X111Y116_ALUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLL_R_X73Y116_SLICE_X111Y116_AO5),
.O6(CLBLL_R_X73Y116_SLICE_X111Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y116_SLICE_X111Y116_MUXF7A (
.I0(CLBLL_R_X73Y116_SLICE_X111Y116_BO6),
.I1(CLBLL_R_X73Y116_SLICE_X111Y116_AO6),
.O(CLBLL_R_X73Y116_SLICE_X111Y116_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y116_SLICE_X111Y116_MUXF7B (
.I0(CLBLL_R_X73Y116_SLICE_X111Y116_DO6),
.I1(CLBLL_R_X73Y116_SLICE_X111Y116_CO6),
.O(CLBLL_R_X73Y116_SLICE_X111Y116_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y116_SLICE_X111Y116_MUXF8 (
.I0(CLBLL_R_X73Y116_SLICE_X111Y116_F7BMUX_O),
.I1(CLBLL_R_X73Y116_SLICE_X111Y116_F7AMUX_O),
.O(CLBLL_R_X73Y116_SLICE_X111Y116_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcafa00c0cafa0)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_DLUT (
.I0(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.O5(CLBLL_R_X73Y118_SLICE_X110Y118_DO5),
.O6(CLBLL_R_X73Y118_SLICE_X110Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddf5a08888f5a0)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.O5(CLBLL_R_X73Y118_SLICE_X110Y118_CO5),
.O6(CLBLL_R_X73Y118_SLICE_X110Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdb97531eca86420)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLL_R_X73Y118_SLICE_X110Y118_BO5),
.O6(CLBLL_R_X73Y118_SLICE_X110Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd75ec64b931a820)
  ) CLBLL_R_X73Y118_SLICE_X110Y118_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.O5(CLBLL_R_X73Y118_SLICE_X110Y118_AO5),
.O6(CLBLL_R_X73Y118_SLICE_X110Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y118_SLICE_X110Y118_MUXF7A (
.I0(CLBLL_R_X73Y118_SLICE_X110Y118_BO6),
.I1(CLBLL_R_X73Y118_SLICE_X110Y118_AO6),
.O(CLBLL_R_X73Y118_SLICE_X110Y118_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y118_SLICE_X110Y118_MUXF7B (
.I0(CLBLL_R_X73Y118_SLICE_X110Y118_DO6),
.I1(CLBLL_R_X73Y118_SLICE_X110Y118_CO6),
.O(CLBLL_R_X73Y118_SLICE_X110Y118_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y118_SLICE_X110Y118_MUXF8 (
.I0(CLBLL_R_X73Y118_SLICE_X110Y118_F7BMUX_O),
.I1(CLBLL_R_X73Y118_SLICE_X110Y118_F7AMUX_O),
.O(CLBLL_R_X73Y118_SLICE_X110Y118_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y118_SLICE_X111Y118_DO5),
.O6(CLBLL_R_X73Y118_SLICE_X111Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y118_SLICE_X111Y118_CO5),
.O6(CLBLL_R_X73Y118_SLICE_X111Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaa00aa)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_BLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y118_SLICE_X111Y118_BO5),
.O6(CLBLL_R_X73Y118_SLICE_X111Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef4aea45e540e04)
  ) CLBLL_R_X73Y118_SLICE_X111Y118_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.O5(CLBLL_R_X73Y118_SLICE_X111Y118_AO5),
.O6(CLBLL_R_X73Y118_SLICE_X111Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y118_SLICE_X111Y118_MUXF7A (
.I0(CLBLL_R_X73Y118_SLICE_X111Y118_BO6),
.I1(CLBLL_R_X73Y118_SLICE_X111Y118_AO6),
.O(CLBLL_R_X73Y118_SLICE_X111Y118_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hef2fe323ec2ce020)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_DLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.O5(CLBLL_R_X73Y119_SLICE_X110Y119_DO5),
.O6(CLBLL_R_X73Y119_SLICE_X110Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef4fe545ea4ae040)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_CLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I4(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.O5(CLBLL_R_X73Y119_SLICE_X110Y119_CO5),
.O6(CLBLL_R_X73Y119_SLICE_X110Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcce2e23300e2e2)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_BLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLL_R_X73Y119_SLICE_X110Y119_BO5),
.O6(CLBLL_R_X73Y119_SLICE_X110Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb833b8ccb800b8)
  ) CLBLL_R_X73Y119_SLICE_X110Y119_ALUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.O5(CLBLL_R_X73Y119_SLICE_X110Y119_AO5),
.O6(CLBLL_R_X73Y119_SLICE_X110Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y119_SLICE_X110Y119_MUXF7A (
.I0(CLBLL_R_X73Y119_SLICE_X110Y119_BO6),
.I1(CLBLL_R_X73Y119_SLICE_X110Y119_AO6),
.O(CLBLL_R_X73Y119_SLICE_X110Y119_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y119_SLICE_X110Y119_MUXF7B (
.I0(CLBLL_R_X73Y119_SLICE_X110Y119_DO6),
.I1(CLBLL_R_X73Y119_SLICE_X110Y119_CO6),
.O(CLBLL_R_X73Y119_SLICE_X110Y119_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y119_SLICE_X110Y119_MUXF8 (
.I0(CLBLL_R_X73Y119_SLICE_X110Y119_F7BMUX_O),
.I1(CLBLL_R_X73Y119_SLICE_X110Y119_F7AMUX_O),
.O(CLBLL_R_X73Y119_SLICE_X110Y119_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa6666aaaa6666)
  ) CLBLL_R_X73Y119_SLICE_X111Y119_DLUT (
.I0(LIOB33_X0Y85_IOB_X0Y85_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(1'b1),
.O5(CLBLL_R_X73Y119_SLICE_X111Y119_DO5),
.O6(CLBLL_R_X73Y119_SLICE_X111Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h556595a55a6a9aaa)
  ) CLBLL_R_X73Y119_SLICE_X111Y119_CLUT (
.I0(CLBLM_L_X70Y123_SLICE_X105Y123_CO6),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_F7AMUX_O),
.I4(CLBLL_R_X73Y118_SLICE_X111Y118_F7AMUX_O),
.I5(CLBLM_L_X74Y119_SLICE_X112Y119_F8MUX_O),
.O5(CLBLL_R_X73Y119_SLICE_X111Y119_CO5),
.O6(CLBLL_R_X73Y119_SLICE_X111Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe4aae455e400e4)
  ) CLBLL_R_X73Y119_SLICE_X111Y119_BLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I5(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.O5(CLBLL_R_X73Y119_SLICE_X111Y119_BO5),
.O6(CLBLL_R_X73Y119_SLICE_X111Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ddddfa508888)
  ) CLBLL_R_X73Y119_SLICE_X111Y119_ALUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.O5(CLBLL_R_X73Y119_SLICE_X111Y119_AO5),
.O6(CLBLL_R_X73Y119_SLICE_X111Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y119_SLICE_X111Y119_MUXF7A (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_BO6),
.I1(CLBLL_R_X73Y119_SLICE_X111Y119_AO6),
.O(CLBLL_R_X73Y119_SLICE_X111Y119_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00aaaaf0f0)
  ) CLBLL_R_X73Y120_SLICE_X110Y120_DLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y120_SLICE_X110Y120_DO5),
.O6(CLBLL_R_X73Y120_SLICE_X110Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdad5d0df8a85808)
  ) CLBLL_R_X73Y120_SLICE_X110Y120_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.O5(CLBLL_R_X73Y120_SLICE_X110Y120_CO5),
.O6(CLBLL_R_X73Y120_SLICE_X110Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heef5eea044f544a0)
  ) CLBLL_R_X73Y120_SLICE_X110Y120_BLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I2(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.O5(CLBLL_R_X73Y120_SLICE_X110Y120_BO5),
.O6(CLBLL_R_X73Y120_SLICE_X110Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5ee44a0a0ee44)
  ) CLBLL_R_X73Y120_SLICE_X110Y120_ALUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.O5(CLBLL_R_X73Y120_SLICE_X110Y120_AO5),
.O6(CLBLL_R_X73Y120_SLICE_X110Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y120_SLICE_X110Y120_MUXF7A (
.I0(CLBLL_R_X73Y120_SLICE_X110Y120_BO6),
.I1(CLBLL_R_X73Y120_SLICE_X110Y120_AO6),
.O(CLBLL_R_X73Y120_SLICE_X110Y120_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y120_SLICE_X110Y120_MUXF7B (
.I0(CLBLL_R_X73Y120_SLICE_X110Y120_DO6),
.I1(CLBLL_R_X73Y120_SLICE_X110Y120_CO6),
.O(CLBLL_R_X73Y120_SLICE_X110Y120_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1eb41eb40f0ff0f0)
  ) CLBLL_R_X73Y120_SLICE_X111Y120_DLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(CLBLL_R_X73Y121_SLICE_X111Y121_F7AMUX_O),
.I2(CLBLM_L_X70Y123_SLICE_X105Y123_CO6),
.I3(CLBLL_R_X73Y120_SLICE_X111Y120_F7AMUX_O),
.I4(CLBLM_L_X74Y120_SLICE_X112Y120_F8MUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLL_R_X73Y120_SLICE_X111Y120_DO5),
.O6(CLBLL_R_X73Y120_SLICE_X111Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11bbee440f0ff0f0)
  ) CLBLL_R_X73Y120_SLICE_X111Y120_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(CLBLL_R_X73Y120_SLICE_X110Y120_F7AMUX_O),
.I2(CLBLL_R_X75Y120_SLICE_X114Y120_F8MUX_O),
.I3(CLBLL_R_X73Y120_SLICE_X110Y120_F7BMUX_O),
.I4(CLBLL_R_X71Y131_SLICE_X107Y131_DO6),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLL_R_X73Y120_SLICE_X111Y120_CO5),
.O6(CLBLL_R_X73Y120_SLICE_X111Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbf3bbc088f388c0)
  ) CLBLL_R_X73Y120_SLICE_X111Y120_BLUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLL_R_X73Y120_SLICE_X111Y120_BO5),
.O6(CLBLL_R_X73Y120_SLICE_X111Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0fff000)
  ) CLBLL_R_X73Y120_SLICE_X111Y120_ALUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I2(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLL_R_X73Y120_SLICE_X111Y120_AO5),
.O6(CLBLL_R_X73Y120_SLICE_X111Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y120_SLICE_X111Y120_MUXF7A (
.I0(CLBLL_R_X73Y120_SLICE_X111Y120_BO6),
.I1(CLBLL_R_X73Y120_SLICE_X111Y120_AO6),
.O(CLBLL_R_X73Y120_SLICE_X111Y120_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y121_SLICE_X110Y121_DO5),
.O6(CLBLL_R_X73Y121_SLICE_X110Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa5a5a66665a5a)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_CLUT (
.I0(CLBLM_L_X70Y129_SLICE_X104Y129_CO6),
.I1(CLBLL_R_X73Y121_SLICE_X111Y121_F7BMUX_O),
.I2(CLBLM_L_X74Y121_SLICE_X112Y121_F8MUX_O),
.I3(CLBLL_R_X73Y121_SLICE_X110Y121_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X73Y121_SLICE_X110Y121_CO5),
.O6(CLBLL_R_X73Y121_SLICE_X110Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfc88fcbb308830)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_BLUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.O5(CLBLL_R_X73Y121_SLICE_X110Y121_BO5),
.O6(CLBLL_R_X73Y121_SLICE_X110Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaae4e45500e4e4)
  ) CLBLL_R_X73Y121_SLICE_X110Y121_ALUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I3(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.O5(CLBLL_R_X73Y121_SLICE_X110Y121_AO5),
.O6(CLBLL_R_X73Y121_SLICE_X110Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y121_SLICE_X110Y121_MUXF7A (
.I0(CLBLL_R_X73Y121_SLICE_X110Y121_BO6),
.I1(CLBLL_R_X73Y121_SLICE_X110Y121_AO6),
.O(CLBLL_R_X73Y121_SLICE_X110Y121_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55e4e4aa00e4e4)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.O5(CLBLL_R_X73Y121_SLICE_X111Y121_DO5),
.O6(CLBLL_R_X73Y121_SLICE_X111Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ffaaccf000aa)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_CLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I1(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.O5(CLBLL_R_X73Y121_SLICE_X111Y121_CO5),
.O6(CLBLL_R_X73Y121_SLICE_X111Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe54f45eae04a40)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_BLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I4(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.O5(CLBLL_R_X73Y121_SLICE_X111Y121_BO5),
.O6(CLBLL_R_X73Y121_SLICE_X111Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeae5e04f4a4540)
  ) CLBLL_R_X73Y121_SLICE_X111Y121_ALUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.O5(CLBLL_R_X73Y121_SLICE_X111Y121_AO5),
.O6(CLBLL_R_X73Y121_SLICE_X111Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y121_SLICE_X111Y121_MUXF7A (
.I0(CLBLL_R_X73Y121_SLICE_X111Y121_BO6),
.I1(CLBLL_R_X73Y121_SLICE_X111Y121_AO6),
.O(CLBLL_R_X73Y121_SLICE_X111Y121_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y121_SLICE_X111Y121_MUXF7B (
.I0(CLBLL_R_X73Y121_SLICE_X111Y121_DO6),
.I1(CLBLL_R_X73Y121_SLICE_X111Y121_CO6),
.O(CLBLL_R_X73Y121_SLICE_X111Y121_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2b5a6492d4656b9)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_DLUT (
.I0(CLBLM_L_X74Y125_SLICE_X112Y125_DO6),
.I1(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I2(CLBLL_R_X73Y123_SLICE_X110Y123_DO6),
.I3(CLBLM_L_X74Y123_SLICE_X112Y123_CO6),
.I4(CLBLL_R_X73Y123_SLICE_X110Y123_CO6),
.I5(CLBLM_L_X72Y122_SLICE_X108Y122_AO6),
.O5(CLBLL_R_X73Y122_SLICE_X110Y122_DO5),
.O6(CLBLL_R_X73Y122_SLICE_X110Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h709fdb24cb1414eb)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_CLUT (
.I0(CLBLM_L_X74Y125_SLICE_X112Y125_DO6),
.I1(CLBLM_L_X74Y123_SLICE_X112Y123_CO6),
.I2(CLBLL_R_X73Y123_SLICE_X110Y123_DO6),
.I3(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.I4(CLBLL_R_X73Y123_SLICE_X110Y123_CO6),
.I5(CLBLM_L_X72Y122_SLICE_X108Y122_AO6),
.O5(CLBLL_R_X73Y122_SLICE_X110Y122_CO5),
.O6(CLBLL_R_X73Y122_SLICE_X110Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a593da46975c619)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_BLUT (
.I0(CLBLL_R_X73Y123_SLICE_X110Y123_DO6),
.I1(CLBLL_R_X73Y123_SLICE_X110Y123_CO6),
.I2(CLBLM_L_X74Y123_SLICE_X112Y123_CO6),
.I3(CLBLM_L_X72Y122_SLICE_X108Y122_AO6),
.I4(CLBLM_L_X74Y125_SLICE_X112Y125_DO6),
.I5(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.O5(CLBLL_R_X73Y122_SLICE_X110Y122_BO5),
.O6(CLBLL_R_X73Y122_SLICE_X110Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h86d3d5a2a695384f)
  ) CLBLL_R_X73Y122_SLICE_X110Y122_ALUT (
.I0(CLBLL_R_X73Y123_SLICE_X110Y123_DO6),
.I1(CLBLL_R_X73Y123_SLICE_X110Y123_CO6),
.I2(CLBLM_L_X74Y125_SLICE_X112Y125_DO6),
.I3(CLBLM_L_X72Y122_SLICE_X108Y122_AO6),
.I4(CLBLM_L_X74Y123_SLICE_X112Y123_CO6),
.I5(CLBLL_R_X75Y123_SLICE_X114Y123_AO6),
.O5(CLBLL_R_X73Y122_SLICE_X110Y122_AO5),
.O6(CLBLL_R_X73Y122_SLICE_X110Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y122_SLICE_X111Y122_DO5),
.O6(CLBLL_R_X73Y122_SLICE_X111Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y122_SLICE_X111Y122_CO5),
.O6(CLBLL_R_X73Y122_SLICE_X111Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y122_SLICE_X111Y122_BO5),
.O6(CLBLL_R_X73Y122_SLICE_X111Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y122_SLICE_X111Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y122_SLICE_X111Y122_AO5),
.O6(CLBLL_R_X73Y122_SLICE_X111Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05af2727fa50d8d8)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_DLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLL_R_X73Y124_SLICE_X111Y124_F7AMUX_O),
.I2(CLBLM_L_X74Y124_SLICE_X112Y124_F8MUX_O),
.I3(CLBLL_R_X73Y124_SLICE_X111Y124_F7BMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.O5(CLBLL_R_X73Y123_SLICE_X110Y123_DO5),
.O6(CLBLL_R_X73Y123_SLICE_X110Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h272705afd8d8fa50)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X74Y123_SLICE_X112Y123_F7AMUX_O),
.I2(CLBLL_R_X73Y123_SLICE_X111Y123_F8MUX_O),
.I3(CLBLL_R_X73Y123_SLICE_X110Y123_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_L_X2Y118_SLICE_X0Y118_CO6),
.O5(CLBLL_R_X73Y123_SLICE_X110Y123_CO5),
.O6(CLBLL_R_X73Y123_SLICE_X110Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe76ba32dc549810)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I3(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.O5(CLBLL_R_X73Y123_SLICE_X110Y123_BO5),
.O6(CLBLL_R_X73Y123_SLICE_X110Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe2cce233e200e2)
  ) CLBLL_R_X73Y123_SLICE_X110Y123_ALUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.O5(CLBLL_R_X73Y123_SLICE_X110Y123_AO5),
.O6(CLBLL_R_X73Y123_SLICE_X110Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y123_SLICE_X110Y123_MUXF7A (
.I0(CLBLL_R_X73Y123_SLICE_X110Y123_BO6),
.I1(CLBLL_R_X73Y123_SLICE_X110Y123_AO6),
.O(CLBLL_R_X73Y123_SLICE_X110Y123_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000acacacac)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_DLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I4(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X73Y123_SLICE_X111Y123_DO5),
.O6(CLBLL_R_X73Y123_SLICE_X111Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50dddd8888)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I2(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X73Y123_SLICE_X111Y123_CO5),
.O6(CLBLL_R_X73Y123_SLICE_X111Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafff0ccaa00f0cc)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_BLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I2(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.O5(CLBLL_R_X73Y123_SLICE_X111Y123_BO5),
.O6(CLBLL_R_X73Y123_SLICE_X111Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44ee44)
  ) CLBLL_R_X73Y123_SLICE_X111Y123_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I3(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I4(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X73Y123_SLICE_X111Y123_AO5),
.O6(CLBLL_R_X73Y123_SLICE_X111Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y123_SLICE_X111Y123_MUXF7A (
.I0(CLBLL_R_X73Y123_SLICE_X111Y123_BO6),
.I1(CLBLL_R_X73Y123_SLICE_X111Y123_AO6),
.O(CLBLL_R_X73Y123_SLICE_X111Y123_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y123_SLICE_X111Y123_MUXF7B (
.I0(CLBLL_R_X73Y123_SLICE_X111Y123_DO6),
.I1(CLBLL_R_X73Y123_SLICE_X111Y123_CO6),
.O(CLBLL_R_X73Y123_SLICE_X111Y123_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y123_SLICE_X111Y123_MUXF8 (
.I0(CLBLL_R_X73Y123_SLICE_X111Y123_F7BMUX_O),
.I1(CLBLL_R_X73Y123_SLICE_X111Y123_F7AMUX_O),
.O(CLBLL_R_X73Y123_SLICE_X111Y123_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcaf0caffca00ca0)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_DLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.O5(CLBLL_R_X73Y124_SLICE_X110Y124_DO5),
.O6(CLBLL_R_X73Y124_SLICE_X110Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffacf0ac0fac00ac)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_CLUT (
.I0(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I1(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.O5(CLBLL_R_X73Y124_SLICE_X110Y124_CO5),
.O6(CLBLL_R_X73Y124_SLICE_X110Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb3bf838cb0bc808)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_BLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I5(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.O5(CLBLL_R_X73Y124_SLICE_X110Y124_BO5),
.O6(CLBLL_R_X73Y124_SLICE_X110Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafcfafc0a0cfa0c0)
  ) CLBLL_R_X73Y124_SLICE_X110Y124_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.O5(CLBLL_R_X73Y124_SLICE_X110Y124_AO5),
.O6(CLBLL_R_X73Y124_SLICE_X110Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y124_SLICE_X110Y124_MUXF7A (
.I0(CLBLL_R_X73Y124_SLICE_X110Y124_BO6),
.I1(CLBLL_R_X73Y124_SLICE_X110Y124_AO6),
.O(CLBLL_R_X73Y124_SLICE_X110Y124_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y124_SLICE_X110Y124_MUXF7B (
.I0(CLBLL_R_X73Y124_SLICE_X110Y124_DO6),
.I1(CLBLL_R_X73Y124_SLICE_X110Y124_CO6),
.O(CLBLL_R_X73Y124_SLICE_X110Y124_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y124_SLICE_X110Y124_MUXF8 (
.I0(CLBLL_R_X73Y124_SLICE_X110Y124_F7BMUX_O),
.I1(CLBLL_R_X73Y124_SLICE_X110Y124_F7AMUX_O),
.O(CLBLL_R_X73Y124_SLICE_X110Y124_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacffacf0ac0fac00)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_DLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.O5(CLBLL_R_X73Y124_SLICE_X111Y124_DO5),
.O6(CLBLL_R_X73Y124_SLICE_X111Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0aaf0aa)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_CLUT (
.I0(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I1(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y124_SLICE_X111Y124_CO5),
.O6(CLBLL_R_X73Y124_SLICE_X111Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_BLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X73Y124_SLICE_X111Y124_BO5),
.O6(CLBLL_R_X73Y124_SLICE_X111Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fcfc0c0c)
  ) CLBLL_R_X73Y124_SLICE_X111Y124_ALUT (
.I0(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I4(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X73Y124_SLICE_X111Y124_AO5),
.O6(CLBLL_R_X73Y124_SLICE_X111Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y124_SLICE_X111Y124_MUXF7A (
.I0(CLBLL_R_X73Y124_SLICE_X111Y124_BO6),
.I1(CLBLL_R_X73Y124_SLICE_X111Y124_AO6),
.O(CLBLL_R_X73Y124_SLICE_X111Y124_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y124_SLICE_X111Y124_MUXF7B (
.I0(CLBLL_R_X73Y124_SLICE_X111Y124_DO6),
.I1(CLBLL_R_X73Y124_SLICE_X111Y124_CO6),
.O(CLBLL_R_X73Y124_SLICE_X111Y124_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ccccaaaa)
  ) CLBLL_R_X73Y125_SLICE_X110Y125_DLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I3(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X73Y125_SLICE_X110Y125_DO5),
.O6(CLBLL_R_X73Y125_SLICE_X110Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ffd8aad855d800)
  ) CLBLL_R_X73Y125_SLICE_X110Y125_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.O5(CLBLL_R_X73Y125_SLICE_X110Y125_CO5),
.O6(CLBLL_R_X73Y125_SLICE_X110Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ccaaccaa)
  ) CLBLL_R_X73Y125_SLICE_X110Y125_BLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I1(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X73Y125_SLICE_X110Y125_BO5),
.O6(CLBLL_R_X73Y125_SLICE_X110Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeef5a04444f5a0)
  ) CLBLL_R_X73Y125_SLICE_X110Y125_ALUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I2(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.O5(CLBLL_R_X73Y125_SLICE_X110Y125_AO5),
.O6(CLBLL_R_X73Y125_SLICE_X110Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y125_SLICE_X110Y125_MUXF7A (
.I0(CLBLL_R_X73Y125_SLICE_X110Y125_BO6),
.I1(CLBLL_R_X73Y125_SLICE_X110Y125_AO6),
.O(CLBLL_R_X73Y125_SLICE_X110Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y125_SLICE_X110Y125_MUXF7B (
.I0(CLBLL_R_X73Y125_SLICE_X110Y125_DO6),
.I1(CLBLL_R_X73Y125_SLICE_X110Y125_CO6),
.O(CLBLL_R_X73Y125_SLICE_X110Y125_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y125_SLICE_X110Y125_MUXF8 (
.I0(CLBLL_R_X73Y125_SLICE_X110Y125_F7BMUX_O),
.I1(CLBLL_R_X73Y125_SLICE_X110Y125_F7AMUX_O),
.O(CLBLL_R_X73Y125_SLICE_X110Y125_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0afafa0a0)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_DLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I1(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I4(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y125_SLICE_X111Y125_DO5),
.O6(CLBLL_R_X73Y125_SLICE_X111Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22f3f3ee22c0c0)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_CLUT (
.I0(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.O5(CLBLL_R_X73Y125_SLICE_X111Y125_CO5),
.O6(CLBLL_R_X73Y125_SLICE_X111Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfebadc9876325410)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I5(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.O5(CLBLL_R_X73Y125_SLICE_X111Y125_BO5),
.O6(CLBLL_R_X73Y125_SLICE_X111Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefc302222fc30)
  ) CLBLL_R_X73Y125_SLICE_X111Y125_ALUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.O5(CLBLL_R_X73Y125_SLICE_X111Y125_AO5),
.O6(CLBLL_R_X73Y125_SLICE_X111Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y125_SLICE_X111Y125_MUXF7A (
.I0(CLBLL_R_X73Y125_SLICE_X111Y125_BO6),
.I1(CLBLL_R_X73Y125_SLICE_X111Y125_AO6),
.O(CLBLL_R_X73Y125_SLICE_X111Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y125_SLICE_X111Y125_MUXF7B (
.I0(CLBLL_R_X73Y125_SLICE_X111Y125_DO6),
.I1(CLBLL_R_X73Y125_SLICE_X111Y125_CO6),
.O(CLBLL_R_X73Y125_SLICE_X111Y125_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y125_SLICE_X111Y125_MUXF8 (
.I0(CLBLL_R_X73Y125_SLICE_X111Y125_F7BMUX_O),
.I1(CLBLL_R_X73Y125_SLICE_X111Y125_F7AMUX_O),
.O(CLBLL_R_X73Y125_SLICE_X111Y125_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbea7362d9c85140)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_DLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.O5(CLBLL_R_X73Y126_SLICE_X110Y126_DO5),
.O6(CLBLL_R_X73Y126_SLICE_X110Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaae4e45500e4e4)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.O5(CLBLL_R_X73Y126_SLICE_X110Y126_CO5),
.O6(CLBLL_R_X73Y126_SLICE_X110Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaaaff00)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_BLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y126_SLICE_X110Y126_BO5),
.O6(CLBLL_R_X73Y126_SLICE_X110Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ddddfa508888)
  ) CLBLL_R_X73Y126_SLICE_X110Y126_ALUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.O5(CLBLL_R_X73Y126_SLICE_X110Y126_AO5),
.O6(CLBLL_R_X73Y126_SLICE_X110Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y126_SLICE_X110Y126_MUXF7A (
.I0(CLBLL_R_X73Y126_SLICE_X110Y126_BO6),
.I1(CLBLL_R_X73Y126_SLICE_X110Y126_AO6),
.O(CLBLL_R_X73Y126_SLICE_X110Y126_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y126_SLICE_X110Y126_MUXF7B (
.I0(CLBLL_R_X73Y126_SLICE_X110Y126_DO6),
.I1(CLBLL_R_X73Y126_SLICE_X110Y126_CO6),
.O(CLBLL_R_X73Y126_SLICE_X110Y126_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y126_SLICE_X110Y126_MUXF8 (
.I0(CLBLL_R_X73Y126_SLICE_X110Y126_F7BMUX_O),
.I1(CLBLL_R_X73Y126_SLICE_X110Y126_F7AMUX_O),
.O(CLBLL_R_X73Y126_SLICE_X110Y126_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4ff55e4e4aa00)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_DLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I2(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.O5(CLBLL_R_X73Y126_SLICE_X111Y126_DO5),
.O6(CLBLL_R_X73Y126_SLICE_X111Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcffacf0ac0fac00a)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_CLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.O5(CLBLL_R_X73Y126_SLICE_X111Y126_CO5),
.O6(CLBLL_R_X73Y126_SLICE_X111Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4ff55e4e4aa00)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.O5(CLBLL_R_X73Y126_SLICE_X111Y126_BO5),
.O6(CLBLL_R_X73Y126_SLICE_X111Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacffacf0ac0fac00)
  ) CLBLL_R_X73Y126_SLICE_X111Y126_ALUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.O5(CLBLL_R_X73Y126_SLICE_X111Y126_AO5),
.O6(CLBLL_R_X73Y126_SLICE_X111Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y126_SLICE_X111Y126_MUXF7A (
.I0(CLBLL_R_X73Y126_SLICE_X111Y126_BO6),
.I1(CLBLL_R_X73Y126_SLICE_X111Y126_AO6),
.O(CLBLL_R_X73Y126_SLICE_X111Y126_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y126_SLICE_X111Y126_MUXF7B (
.I0(CLBLL_R_X73Y126_SLICE_X111Y126_DO6),
.I1(CLBLL_R_X73Y126_SLICE_X111Y126_CO6),
.O(CLBLL_R_X73Y126_SLICE_X111Y126_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heef5eea044f544a0)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_DLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I2(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.O5(CLBLL_R_X73Y127_SLICE_X110Y127_DO5),
.O6(CLBLL_R_X73Y127_SLICE_X110Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd5df858ad0da808)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_CLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I4(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.O5(CLBLL_R_X73Y127_SLICE_X110Y127_CO5),
.O6(CLBLL_R_X73Y127_SLICE_X110Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeefa504444fa50)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.O5(CLBLL_R_X73Y127_SLICE_X110Y127_BO5),
.O6(CLBLL_R_X73Y127_SLICE_X110Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ccaa00f0ccaa)
  ) CLBLL_R_X73Y127_SLICE_X110Y127_ALUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I1(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I2(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.O5(CLBLL_R_X73Y127_SLICE_X110Y127_AO5),
.O6(CLBLL_R_X73Y127_SLICE_X110Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y127_SLICE_X110Y127_MUXF7A (
.I0(CLBLL_R_X73Y127_SLICE_X110Y127_BO6),
.I1(CLBLL_R_X73Y127_SLICE_X110Y127_AO6),
.O(CLBLL_R_X73Y127_SLICE_X110Y127_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y127_SLICE_X110Y127_MUXF7B (
.I0(CLBLL_R_X73Y127_SLICE_X110Y127_DO6),
.I1(CLBLL_R_X73Y127_SLICE_X110Y127_CO6),
.O(CLBLL_R_X73Y127_SLICE_X110Y127_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y127_SLICE_X110Y127_MUXF8 (
.I0(CLBLL_R_X73Y127_SLICE_X110Y127_F7BMUX_O),
.I1(CLBLL_R_X73Y127_SLICE_X110Y127_F7AMUX_O),
.O(CLBLL_R_X73Y127_SLICE_X110Y127_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y127_SLICE_X111Y127_DO5),
.O6(CLBLL_R_X73Y127_SLICE_X111Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa5a5a66665a5a)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_CLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.I1(CLBLM_L_X74Y127_SLICE_X112Y127_F7AMUX_O),
.I2(CLBLL_R_X73Y127_SLICE_X110Y127_F8MUX_O),
.I3(CLBLL_R_X73Y127_SLICE_X111Y127_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X73Y127_SLICE_X111Y127_CO5),
.O6(CLBLL_R_X73Y127_SLICE_X111Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf8fda8ad585d080)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I4(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.O5(CLBLL_R_X73Y127_SLICE_X111Y127_BO5),
.O6(CLBLL_R_X73Y127_SLICE_X111Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afcfcfa0a0c0c)
  ) CLBLL_R_X73Y127_SLICE_X111Y127_ALUT (
.I0(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.O5(CLBLL_R_X73Y127_SLICE_X111Y127_AO5),
.O6(CLBLL_R_X73Y127_SLICE_X111Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y127_SLICE_X111Y127_MUXF7A (
.I0(CLBLL_R_X73Y127_SLICE_X111Y127_BO6),
.I1(CLBLL_R_X73Y127_SLICE_X111Y127_AO6),
.O(CLBLL_R_X73Y127_SLICE_X111Y127_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44ee44)
  ) CLBLL_R_X73Y128_SLICE_X110Y128_DLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y128_SLICE_X110Y128_DO5),
.O6(CLBLL_R_X73Y128_SLICE_X110Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00aaaaf0f0)
  ) CLBLL_R_X73Y128_SLICE_X110Y128_CLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X73Y128_SLICE_X110Y128_CO5),
.O6(CLBLL_R_X73Y128_SLICE_X110Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfd58f85dad08a80)
  ) CLBLL_R_X73Y128_SLICE_X110Y128_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I5(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.O5(CLBLL_R_X73Y128_SLICE_X110Y128_BO5),
.O6(CLBLL_R_X73Y128_SLICE_X110Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe5eae04f454a40)
  ) CLBLL_R_X73Y128_SLICE_X110Y128_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.O5(CLBLL_R_X73Y128_SLICE_X110Y128_AO5),
.O6(CLBLL_R_X73Y128_SLICE_X110Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y128_SLICE_X110Y128_MUXF7A (
.I0(CLBLL_R_X73Y128_SLICE_X110Y128_BO6),
.I1(CLBLL_R_X73Y128_SLICE_X110Y128_AO6),
.O(CLBLL_R_X73Y128_SLICE_X110Y128_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y128_SLICE_X110Y128_MUXF7B (
.I0(CLBLL_R_X73Y128_SLICE_X110Y128_DO6),
.I1(CLBLL_R_X73Y128_SLICE_X110Y128_CO6),
.O(CLBLL_R_X73Y128_SLICE_X110Y128_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y128_SLICE_X110Y128_MUXF8 (
.I0(CLBLL_R_X73Y128_SLICE_X110Y128_F7BMUX_O),
.I1(CLBLL_R_X73Y128_SLICE_X110Y128_F7AMUX_O),
.O(CLBLL_R_X73Y128_SLICE_X110Y128_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf8fb383bc8cb080)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_DLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I4(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.O5(CLBLL_R_X73Y128_SLICE_X111Y128_DO5),
.O6(CLBLL_R_X73Y128_SLICE_X111Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_CLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I3(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y128_SLICE_X111Y128_CO5),
.O6(CLBLL_R_X73Y128_SLICE_X111Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ccaa00f0ccaa)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_BLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.O5(CLBLL_R_X73Y128_SLICE_X111Y128_BO5),
.O6(CLBLL_R_X73Y128_SLICE_X111Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dd88dd88)
  ) CLBLL_R_X73Y128_SLICE_X111Y128_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I2(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X73Y128_SLICE_X111Y128_AO5),
.O6(CLBLL_R_X73Y128_SLICE_X111Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y128_SLICE_X111Y128_MUXF7A (
.I0(CLBLL_R_X73Y128_SLICE_X111Y128_BO6),
.I1(CLBLL_R_X73Y128_SLICE_X111Y128_AO6),
.O(CLBLL_R_X73Y128_SLICE_X111Y128_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y128_SLICE_X111Y128_MUXF7B (
.I0(CLBLL_R_X73Y128_SLICE_X111Y128_DO6),
.I1(CLBLL_R_X73Y128_SLICE_X111Y128_CO6),
.O(CLBLL_R_X73Y128_SLICE_X111Y128_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X73Y129_SLICE_X110Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X73Y129_SLICE_X110Y129_DO5),
.O6(CLBLL_R_X73Y129_SLICE_X110Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2727d8d805affa50)
  ) CLBLL_R_X73Y129_SLICE_X110Y129_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X74Y129_SLICE_X112Y129_F7AMUX_O),
.I2(CLBLL_R_X73Y129_SLICE_X111Y129_F8MUX_O),
.I3(CLBLL_R_X73Y129_SLICE_X110Y129_F7AMUX_O),
.I4(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X73Y129_SLICE_X110Y129_CO5),
.O6(CLBLL_R_X73Y129_SLICE_X110Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22fcfc3030)
  ) CLBLL_R_X73Y129_SLICE_X110Y129_BLUT (
.I0(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y129_SLICE_X110Y129_BO5),
.O6(CLBLL_R_X73Y129_SLICE_X110Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddf5a08888f5a0)
  ) CLBLL_R_X73Y129_SLICE_X110Y129_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.O5(CLBLL_R_X73Y129_SLICE_X110Y129_AO5),
.O6(CLBLL_R_X73Y129_SLICE_X110Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y129_SLICE_X110Y129_MUXF7A (
.I0(CLBLL_R_X73Y129_SLICE_X110Y129_BO6),
.I1(CLBLL_R_X73Y129_SLICE_X110Y129_AO6),
.O(CLBLL_R_X73Y129_SLICE_X110Y129_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cfcfafa0c0c0)
  ) CLBLL_R_X73Y129_SLICE_X111Y129_DLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.O5(CLBLL_R_X73Y129_SLICE_X111Y129_DO5),
.O6(CLBLL_R_X73Y129_SLICE_X111Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeae5e0ef4a45404)
  ) CLBLL_R_X73Y129_SLICE_X111Y129_CLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.O5(CLBLL_R_X73Y129_SLICE_X111Y129_CO5),
.O6(CLBLL_R_X73Y129_SLICE_X111Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcffac0facf0ac00a)
  ) CLBLL_R_X73Y129_SLICE_X111Y129_BLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.O5(CLBLL_R_X73Y129_SLICE_X111Y129_BO5),
.O6(CLBLL_R_X73Y129_SLICE_X111Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0aaccaacc)
  ) CLBLL_R_X73Y129_SLICE_X111Y129_ALUT (
.I0(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X73Y129_SLICE_X111Y129_AO5),
.O6(CLBLL_R_X73Y129_SLICE_X111Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y129_SLICE_X111Y129_MUXF7A (
.I0(CLBLL_R_X73Y129_SLICE_X111Y129_BO6),
.I1(CLBLL_R_X73Y129_SLICE_X111Y129_AO6),
.O(CLBLL_R_X73Y129_SLICE_X111Y129_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X73Y129_SLICE_X111Y129_MUXF7B (
.I0(CLBLL_R_X73Y129_SLICE_X111Y129_DO6),
.I1(CLBLL_R_X73Y129_SLICE_X111Y129_CO6),
.O(CLBLL_R_X73Y129_SLICE_X111Y129_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X73Y129_SLICE_X111Y129_MUXF8 (
.I0(CLBLL_R_X73Y129_SLICE_X111Y129_F7BMUX_O),
.I1(CLBLL_R_X73Y129_SLICE_X111Y129_F7AMUX_O),
.O(CLBLL_R_X73Y129_SLICE_X111Y129_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y115_SLICE_X114Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y115_SLICE_X114Y115_DO5),
.O6(CLBLL_R_X75Y115_SLICE_X114Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y115_SLICE_X114Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y115_SLICE_X114Y115_CO5),
.O6(CLBLL_R_X75Y115_SLICE_X114Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55d8d8aa00d8d8)
  ) CLBLL_R_X75Y115_SLICE_X114Y115_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.O5(CLBLL_R_X75Y115_SLICE_X114Y115_BO5),
.O6(CLBLL_R_X75Y115_SLICE_X114Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLL_R_X75Y115_SLICE_X114Y115_ALUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X75Y115_SLICE_X114Y115_AO5),
.O6(CLBLL_R_X75Y115_SLICE_X114Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y115_SLICE_X114Y115_MUXF7A (
.I0(CLBLL_R_X75Y115_SLICE_X114Y115_BO6),
.I1(CLBLL_R_X75Y115_SLICE_X114Y115_AO6),
.O(CLBLL_R_X75Y115_SLICE_X114Y115_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaafff0ccaa00f0)
  ) CLBLL_R_X75Y115_SLICE_X115Y115_DLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.O5(CLBLL_R_X75Y115_SLICE_X115Y115_DO5),
.O6(CLBLL_R_X75Y115_SLICE_X115Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0eeeef5a04444)
  ) CLBLL_R_X75Y115_SLICE_X115Y115_CLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.O5(CLBLL_R_X75Y115_SLICE_X115Y115_CO5),
.O6(CLBLL_R_X75Y115_SLICE_X115Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ff33cc00)
  ) CLBLL_R_X75Y115_SLICE_X115Y115_BLUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I4(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X75Y115_SLICE_X115Y115_BO5),
.O6(CLBLL_R_X75Y115_SLICE_X115Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7d5e6c4b391a280)
  ) CLBLL_R_X75Y115_SLICE_X115Y115_ALUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I3(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.O5(CLBLL_R_X75Y115_SLICE_X115Y115_AO5),
.O6(CLBLL_R_X75Y115_SLICE_X115Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y115_SLICE_X115Y115_MUXF7A (
.I0(CLBLL_R_X75Y115_SLICE_X115Y115_BO6),
.I1(CLBLL_R_X75Y115_SLICE_X115Y115_AO6),
.O(CLBLL_R_X75Y115_SLICE_X115Y115_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y115_SLICE_X115Y115_MUXF7B (
.I0(CLBLL_R_X75Y115_SLICE_X115Y115_DO6),
.I1(CLBLL_R_X75Y115_SLICE_X115Y115_CO6),
.O(CLBLL_R_X75Y115_SLICE_X115Y115_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X75Y115_SLICE_X115Y115_MUXF8 (
.I0(CLBLL_R_X75Y115_SLICE_X115Y115_F7BMUX_O),
.I1(CLBLL_R_X75Y115_SLICE_X115Y115_F7AMUX_O),
.O(CLBLL_R_X75Y115_SLICE_X115Y115_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y116_SLICE_X114Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y116_SLICE_X114Y116_DO5),
.O6(CLBLL_R_X75Y116_SLICE_X114Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h272705afd8d8fa50)
  ) CLBLL_R_X75Y116_SLICE_X114Y116_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLL_R_X75Y115_SLICE_X114Y115_F7AMUX_O),
.I2(CLBLL_R_X75Y115_SLICE_X115Y115_F8MUX_O),
.I3(CLBLL_R_X75Y116_SLICE_X114Y116_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_R_X71Y131_SLICE_X107Y131_AO6),
.O5(CLBLL_R_X75Y116_SLICE_X114Y116_CO5),
.O6(CLBLL_R_X75Y116_SLICE_X114Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2ffe233e2cce200)
  ) CLBLL_R_X75Y116_SLICE_X114Y116_BLUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.O5(CLBLL_R_X75Y116_SLICE_X114Y116_BO5),
.O6(CLBLL_R_X75Y116_SLICE_X114Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefc22fcee302230)
  ) CLBLL_R_X75Y116_SLICE_X114Y116_ALUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.O5(CLBLL_R_X75Y116_SLICE_X114Y116_AO5),
.O6(CLBLL_R_X75Y116_SLICE_X114Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y116_SLICE_X114Y116_MUXF7A (
.I0(CLBLL_R_X75Y116_SLICE_X114Y116_BO6),
.I1(CLBLL_R_X75Y116_SLICE_X114Y116_AO6),
.O(CLBLL_R_X75Y116_SLICE_X114Y116_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y116_SLICE_X115Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y116_SLICE_X115Y116_DO5),
.O6(CLBLL_R_X75Y116_SLICE_X115Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y116_SLICE_X115Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y116_SLICE_X115Y116_CO5),
.O6(CLBLL_R_X75Y116_SLICE_X115Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfafc0a0cfa0c0a)
  ) CLBLL_R_X75Y116_SLICE_X115Y116_BLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.O5(CLBLL_R_X75Y116_SLICE_X115Y116_BO5),
.O6(CLBLL_R_X75Y116_SLICE_X115Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfacf0acffac00ac0)
  ) CLBLL_R_X75Y116_SLICE_X115Y116_ALUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I5(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.O5(CLBLL_R_X75Y116_SLICE_X115Y116_AO5),
.O6(CLBLL_R_X75Y116_SLICE_X115Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y116_SLICE_X115Y116_MUXF7A (
.I0(CLBLL_R_X75Y116_SLICE_X115Y116_BO6),
.I1(CLBLL_R_X75Y116_SLICE_X115Y116_AO6),
.O(CLBLL_R_X75Y116_SLICE_X115Y116_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8ff55d8d8aa00)
  ) CLBLL_R_X75Y117_SLICE_X114Y117_DLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.O5(CLBLL_R_X75Y117_SLICE_X114Y117_DO5),
.O6(CLBLL_R_X75Y117_SLICE_X114Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5dd88a0a0dd88)
  ) CLBLL_R_X75Y117_SLICE_X114Y117_CLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I3(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.O5(CLBLL_R_X75Y117_SLICE_X114Y117_CO5),
.O6(CLBLL_R_X75Y117_SLICE_X114Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaccccff00)
  ) CLBLL_R_X75Y117_SLICE_X114Y117_BLUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X75Y117_SLICE_X114Y117_BO5),
.O6(CLBLL_R_X75Y117_SLICE_X114Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0aaffccf0aa00)
  ) CLBLL_R_X75Y117_SLICE_X114Y117_ALUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.O5(CLBLL_R_X75Y117_SLICE_X114Y117_AO5),
.O6(CLBLL_R_X75Y117_SLICE_X114Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y117_SLICE_X114Y117_MUXF7A (
.I0(CLBLL_R_X75Y117_SLICE_X114Y117_BO6),
.I1(CLBLL_R_X75Y117_SLICE_X114Y117_AO6),
.O(CLBLL_R_X75Y117_SLICE_X114Y117_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y117_SLICE_X114Y117_MUXF7B (
.I0(CLBLL_R_X75Y117_SLICE_X114Y117_DO6),
.I1(CLBLL_R_X75Y117_SLICE_X114Y117_CO6),
.O(CLBLL_R_X75Y117_SLICE_X114Y117_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00f0f0aaaa)
  ) CLBLL_R_X75Y117_SLICE_X115Y117_DLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X75Y117_SLICE_X115Y117_DO5),
.O6(CLBLL_R_X75Y117_SLICE_X115Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLL_R_X75Y117_SLICE_X115Y117_CLUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X75Y117_SLICE_X115Y117_CO5),
.O6(CLBLL_R_X75Y117_SLICE_X115Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0caca0f00caca)
  ) CLBLL_R_X75Y117_SLICE_X115Y117_BLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.O5(CLBLL_R_X75Y117_SLICE_X115Y117_BO5),
.O6(CLBLL_R_X75Y117_SLICE_X115Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe32f23ece02c20)
  ) CLBLL_R_X75Y117_SLICE_X115Y117_ALUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I5(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.O5(CLBLL_R_X75Y117_SLICE_X115Y117_AO5),
.O6(CLBLL_R_X75Y117_SLICE_X115Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y117_SLICE_X115Y117_MUXF7A (
.I0(CLBLL_R_X75Y117_SLICE_X115Y117_BO6),
.I1(CLBLL_R_X75Y117_SLICE_X115Y117_AO6),
.O(CLBLL_R_X75Y117_SLICE_X115Y117_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y117_SLICE_X115Y117_MUXF7B (
.I0(CLBLL_R_X75Y117_SLICE_X115Y117_DO6),
.I1(CLBLL_R_X75Y117_SLICE_X115Y117_CO6),
.O(CLBLL_R_X75Y117_SLICE_X115Y117_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X75Y117_SLICE_X115Y117_MUXF8 (
.I0(CLBLL_R_X75Y117_SLICE_X115Y117_F7BMUX_O),
.I1(CLBLL_R_X75Y117_SLICE_X115Y117_F7AMUX_O),
.O(CLBLL_R_X75Y117_SLICE_X115Y117_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa55aaaaaa55aa)
  ) CLBLL_R_X75Y118_SLICE_X114Y118_DLUT (
.I0(LIOB33_X0Y85_IOB_X0Y85_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(1'b1),
.O5(CLBLL_R_X75Y118_SLICE_X114Y118_DO5),
.O6(CLBLL_R_X75Y118_SLICE_X114Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05278daffad87250)
  ) CLBLL_R_X75Y118_SLICE_X114Y118_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLL_R_X75Y118_SLICE_X115Y118_F8MUX_O),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_F7AMUX_O),
.I4(CLBLL_R_X75Y119_SLICE_X114Y119_F7AMUX_O),
.I5(CLBLM_L_X70Y128_SLICE_X105Y128_CO6),
.O5(CLBLL_R_X75Y118_SLICE_X114Y118_CO5),
.O6(CLBLL_R_X75Y118_SLICE_X114Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8ff55d8d8aa00)
  ) CLBLL_R_X75Y118_SLICE_X114Y118_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.O5(CLBLL_R_X75Y118_SLICE_X114Y118_BO5),
.O6(CLBLL_R_X75Y118_SLICE_X114Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7b3d591e6a2c480)
  ) CLBLL_R_X75Y118_SLICE_X114Y118_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I5(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.O5(CLBLL_R_X75Y118_SLICE_X114Y118_AO5),
.O6(CLBLL_R_X75Y118_SLICE_X114Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y118_SLICE_X114Y118_MUXF7A (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_BO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_AO6),
.O(CLBLL_R_X75Y118_SLICE_X114Y118_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacafff0caca0f00)
  ) CLBLL_R_X75Y118_SLICE_X115Y118_DLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLL_R_X75Y118_SLICE_X115Y118_DO5),
.O6(CLBLL_R_X75Y118_SLICE_X115Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeae5e04f4a4540)
  ) CLBLL_R_X75Y118_SLICE_X115Y118_CLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I5(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.O5(CLBLL_R_X75Y118_SLICE_X115Y118_CO5),
.O6(CLBLL_R_X75Y118_SLICE_X115Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddfa508888fa50)
  ) CLBLL_R_X75Y118_SLICE_X115Y118_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.O5(CLBLL_R_X75Y118_SLICE_X115Y118_BO5),
.O6(CLBLL_R_X75Y118_SLICE_X115Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeef5a04444f5a0)
  ) CLBLL_R_X75Y118_SLICE_X115Y118_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.O5(CLBLL_R_X75Y118_SLICE_X115Y118_AO5),
.O6(CLBLL_R_X75Y118_SLICE_X115Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y118_SLICE_X115Y118_MUXF7A (
.I0(CLBLL_R_X75Y118_SLICE_X115Y118_BO6),
.I1(CLBLL_R_X75Y118_SLICE_X115Y118_AO6),
.O(CLBLL_R_X75Y118_SLICE_X115Y118_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y118_SLICE_X115Y118_MUXF7B (
.I0(CLBLL_R_X75Y118_SLICE_X115Y118_DO6),
.I1(CLBLL_R_X75Y118_SLICE_X115Y118_CO6),
.O(CLBLL_R_X75Y118_SLICE_X115Y118_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X75Y118_SLICE_X115Y118_MUXF8 (
.I0(CLBLL_R_X75Y118_SLICE_X115Y118_F7BMUX_O),
.I1(CLBLL_R_X75Y118_SLICE_X115Y118_F7AMUX_O),
.O(CLBLL_R_X75Y118_SLICE_X115Y118_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y119_SLICE_X114Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y119_SLICE_X114Y119_DO5),
.O6(CLBLL_R_X75Y119_SLICE_X114Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y119_SLICE_X114Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y119_SLICE_X114Y119_CO5),
.O6(CLBLL_R_X75Y119_SLICE_X114Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee50eefa445044)
  ) CLBLL_R_X75Y119_SLICE_X114Y119_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.O5(CLBLL_R_X75Y119_SLICE_X114Y119_BO5),
.O6(CLBLL_R_X75Y119_SLICE_X114Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hef4fe545ea4ae040)
  ) CLBLL_R_X75Y119_SLICE_X114Y119_ALUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I4(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.O5(CLBLL_R_X75Y119_SLICE_X114Y119_AO5),
.O6(CLBLL_R_X75Y119_SLICE_X114Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y119_SLICE_X114Y119_MUXF7A (
.I0(CLBLL_R_X75Y119_SLICE_X114Y119_BO6),
.I1(CLBLL_R_X75Y119_SLICE_X114Y119_AO6),
.O(CLBLL_R_X75Y119_SLICE_X114Y119_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y119_SLICE_X115Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y119_SLICE_X115Y119_DO5),
.O6(CLBLL_R_X75Y119_SLICE_X115Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y119_SLICE_X115Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y119_SLICE_X115Y119_CO5),
.O6(CLBLL_R_X75Y119_SLICE_X115Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef45e54aea40e04)
  ) CLBLL_R_X75Y119_SLICE_X115Y119_BLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I5(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.O5(CLBLL_R_X75Y119_SLICE_X115Y119_BO5),
.O6(CLBLL_R_X75Y119_SLICE_X115Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe76ba32dc549810)
  ) CLBLL_R_X75Y119_SLICE_X115Y119_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.O5(CLBLL_R_X75Y119_SLICE_X115Y119_AO5),
.O6(CLBLL_R_X75Y119_SLICE_X115Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y119_SLICE_X115Y119_MUXF7A (
.I0(CLBLL_R_X75Y119_SLICE_X115Y119_BO6),
.I1(CLBLL_R_X75Y119_SLICE_X115Y119_AO6),
.O(CLBLL_R_X75Y119_SLICE_X115Y119_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacff0facacf000)
  ) CLBLL_R_X75Y120_SLICE_X114Y120_DLUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.O5(CLBLL_R_X75Y120_SLICE_X114Y120_DO5),
.O6(CLBLL_R_X75Y120_SLICE_X114Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0fcfcafa00c0c)
  ) CLBLL_R_X75Y120_SLICE_X114Y120_CLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.O5(CLBLL_R_X75Y120_SLICE_X114Y120_CO5),
.O6(CLBLL_R_X75Y120_SLICE_X114Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbd9eac873516240)
  ) CLBLL_R_X75Y120_SLICE_X114Y120_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.O5(CLBLL_R_X75Y120_SLICE_X114Y120_BO5),
.O6(CLBLL_R_X75Y120_SLICE_X114Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdb97531eca86420)
  ) CLBLL_R_X75Y120_SLICE_X114Y120_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I2(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.O5(CLBLL_R_X75Y120_SLICE_X114Y120_AO5),
.O6(CLBLL_R_X75Y120_SLICE_X114Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y120_SLICE_X114Y120_MUXF7A (
.I0(CLBLL_R_X75Y120_SLICE_X114Y120_BO6),
.I1(CLBLL_R_X75Y120_SLICE_X114Y120_AO6),
.O(CLBLL_R_X75Y120_SLICE_X114Y120_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y120_SLICE_X114Y120_MUXF7B (
.I0(CLBLL_R_X75Y120_SLICE_X114Y120_DO6),
.I1(CLBLL_R_X75Y120_SLICE_X114Y120_CO6),
.O(CLBLL_R_X75Y120_SLICE_X114Y120_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X75Y120_SLICE_X114Y120_MUXF8 (
.I0(CLBLL_R_X75Y120_SLICE_X114Y120_F7BMUX_O),
.I1(CLBLL_R_X75Y120_SLICE_X114Y120_F7AMUX_O),
.O(CLBLL_R_X75Y120_SLICE_X114Y120_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y120_SLICE_X115Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y120_SLICE_X115Y120_DO5),
.O6(CLBLL_R_X75Y120_SLICE_X115Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55665a5a99aa5a5a)
  ) CLBLL_R_X75Y120_SLICE_X115Y120_CLUT (
.I0(CLBLL_L_X2Y123_SLICE_X0Y123_DO6),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLM_L_X76Y120_SLICE_X116Y120_F8MUX_O),
.I3(CLBLL_R_X75Y120_SLICE_X115Y120_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLL_R_X75Y119_SLICE_X115Y119_F7AMUX_O),
.O5(CLBLL_R_X75Y120_SLICE_X115Y120_CO5),
.O6(CLBLL_R_X75Y120_SLICE_X115Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00e4e4e4e4)
  ) CLBLL_R_X75Y120_SLICE_X115Y120_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I3(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X75Y120_SLICE_X115Y120_BO5),
.O6(CLBLL_R_X75Y120_SLICE_X115Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaccccf0f0)
  ) CLBLL_R_X75Y120_SLICE_X115Y120_ALUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X75Y120_SLICE_X115Y120_AO5),
.O6(CLBLL_R_X75Y120_SLICE_X115Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y120_SLICE_X115Y120_MUXF7A (
.I0(CLBLL_R_X75Y120_SLICE_X115Y120_BO6),
.I1(CLBLL_R_X75Y120_SLICE_X115Y120_AO6),
.O(CLBLL_R_X75Y120_SLICE_X115Y120_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y123_SLICE_X114Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X114Y123_DO5),
.O6(CLBLL_R_X75Y123_SLICE_X114Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y123_SLICE_X114Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X114Y123_CO5),
.O6(CLBLL_R_X75Y123_SLICE_X114Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y123_SLICE_X114Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X114Y123_BO5),
.O6(CLBLL_R_X75Y123_SLICE_X114Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3636c63636c6c6c6)
  ) CLBLL_R_X75Y123_SLICE_X114Y123_ALUT (
.I0(CLBLL_R_X75Y124_SLICE_X114Y124_F8MUX_O),
.I1(CLBLM_L_X70Y121_SLICE_X105Y121_CO6),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(CLBLL_R_X75Y124_SLICE_X115Y124_F7BMUX_O),
.I5(CLBLL_R_X75Y124_SLICE_X115Y124_F7AMUX_O),
.O5(CLBLL_R_X75Y123_SLICE_X114Y123_AO5),
.O6(CLBLL_R_X75Y123_SLICE_X114Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y123_SLICE_X115Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X115Y123_DO5),
.O6(CLBLL_R_X75Y123_SLICE_X115Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y123_SLICE_X115Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X115Y123_CO5),
.O6(CLBLL_R_X75Y123_SLICE_X115Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y123_SLICE_X115Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X115Y123_BO5),
.O6(CLBLL_R_X75Y123_SLICE_X115Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y123_SLICE_X115Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y123_SLICE_X115Y123_AO5),
.O6(CLBLL_R_X75Y123_SLICE_X115Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcee30eefc223022)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_DLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.O5(CLBLL_R_X75Y124_SLICE_X114Y124_DO5),
.O6(CLBLL_R_X75Y124_SLICE_X114Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb3bf838cb0bc808)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_CLUT (
.I0(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.O5(CLBLL_R_X75Y124_SLICE_X114Y124_CO5),
.O6(CLBLL_R_X75Y124_SLICE_X114Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfa0afa0a)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_BLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X75Y124_SLICE_X114Y124_BO5),
.O6(CLBLL_R_X75Y124_SLICE_X114Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbd97351eac86240)
  ) CLBLL_R_X75Y124_SLICE_X114Y124_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I4(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.O5(CLBLL_R_X75Y124_SLICE_X114Y124_AO5),
.O6(CLBLL_R_X75Y124_SLICE_X114Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y124_SLICE_X114Y124_MUXF7A (
.I0(CLBLL_R_X75Y124_SLICE_X114Y124_BO6),
.I1(CLBLL_R_X75Y124_SLICE_X114Y124_AO6),
.O(CLBLL_R_X75Y124_SLICE_X114Y124_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y124_SLICE_X114Y124_MUXF7B (
.I0(CLBLL_R_X75Y124_SLICE_X114Y124_DO6),
.I1(CLBLL_R_X75Y124_SLICE_X114Y124_CO6),
.O(CLBLL_R_X75Y124_SLICE_X114Y124_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X75Y124_SLICE_X114Y124_MUXF8 (
.I0(CLBLL_R_X75Y124_SLICE_X114Y124_F7BMUX_O),
.I1(CLBLL_R_X75Y124_SLICE_X114Y124_F7AMUX_O),
.O(CLBLL_R_X75Y124_SLICE_X114Y124_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffac0facf0ac00ac)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_DLUT (
.I0(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.O5(CLBLL_R_X75Y124_SLICE_X115Y124_DO5),
.O6(CLBLL_R_X75Y124_SLICE_X115Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacffac0facf0ac00)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_CLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I1(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.O5(CLBLL_R_X75Y124_SLICE_X115Y124_CO5),
.O6(CLBLL_R_X75Y124_SLICE_X115Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccf0f0aaaa)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_BLUT (
.I0(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X75Y124_SLICE_X115Y124_BO5),
.O6(CLBLL_R_X75Y124_SLICE_X115Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccf0f0ff00)
  ) CLBLL_R_X75Y124_SLICE_X115Y124_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X75Y124_SLICE_X115Y124_AO5),
.O6(CLBLL_R_X75Y124_SLICE_X115Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y124_SLICE_X115Y124_MUXF7A (
.I0(CLBLL_R_X75Y124_SLICE_X115Y124_BO6),
.I1(CLBLL_R_X75Y124_SLICE_X115Y124_AO6),
.O(CLBLL_R_X75Y124_SLICE_X115Y124_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y124_SLICE_X115Y124_MUXF7B (
.I0(CLBLL_R_X75Y124_SLICE_X115Y124_DO6),
.I1(CLBLL_R_X75Y124_SLICE_X115Y124_CO6),
.O(CLBLL_R_X75Y124_SLICE_X115Y124_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y125_SLICE_X114Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y125_SLICE_X114Y125_DO5),
.O6(CLBLL_R_X75Y125_SLICE_X114Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11bbee440f0ff0f0)
  ) CLBLL_R_X75Y125_SLICE_X114Y125_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(CLBLL_R_X75Y125_SLICE_X115Y125_F7AMUX_O),
.I2(CLBLM_L_X76Y125_SLICE_X116Y125_F8MUX_O),
.I3(CLBLL_R_X75Y125_SLICE_X114Y125_F7AMUX_O),
.I4(CLBLM_L_X70Y121_SLICE_X105Y121_CO6),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLL_R_X75Y125_SLICE_X114Y125_CO5),
.O6(CLBLL_R_X75Y125_SLICE_X114Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLL_R_X75Y125_SLICE_X114Y125_BLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I2(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X75Y125_SLICE_X114Y125_BO5),
.O6(CLBLL_R_X75Y125_SLICE_X114Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888fa50fa50)
  ) CLBLL_R_X75Y125_SLICE_X114Y125_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I2(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I4(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X75Y125_SLICE_X114Y125_AO5),
.O6(CLBLL_R_X75Y125_SLICE_X114Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y125_SLICE_X114Y125_MUXF7A (
.I0(CLBLL_R_X75Y125_SLICE_X114Y125_BO6),
.I1(CLBLL_R_X75Y125_SLICE_X114Y125_AO6),
.O(CLBLL_R_X75Y125_SLICE_X114Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h05faaf5027d827d8)
  ) CLBLL_R_X75Y125_SLICE_X115Y125_DLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X76Y124_SLICE_X116Y124_F7AMUX_O),
.I2(CLBLL_R_X77Y125_SLICE_X118Y125_F8MUX_O),
.I3(CLBLM_L_X70Y122_SLICE_X104Y122_CO6),
.I4(CLBLM_L_X76Y124_SLICE_X116Y124_F7BMUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X75Y125_SLICE_X115Y125_DO5),
.O6(CLBLL_R_X75Y125_SLICE_X115Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4477bb880c3ff3c0)
  ) CLBLL_R_X75Y125_SLICE_X115Y125_CLUT (
.I0(CLBLL_R_X75Y126_SLICE_X115Y126_F7BMUX_O),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(CLBLL_R_X75Y126_SLICE_X115Y126_F7AMUX_O),
.I3(CLBLM_L_X76Y125_SLICE_X117Y125_F8MUX_O),
.I4(CLBLL_R_X71Y131_SLICE_X107Y131_DO6),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X75Y125_SLICE_X115Y125_CO5),
.O6(CLBLL_R_X75Y125_SLICE_X115Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeef3c02222f3c0)
  ) CLBLL_R_X75Y125_SLICE_X115Y125_BLUT (
.I0(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.O5(CLBLL_R_X75Y125_SLICE_X115Y125_BO5),
.O6(CLBLL_R_X75Y125_SLICE_X115Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50dddd8888)
  ) CLBLL_R_X75Y125_SLICE_X115Y125_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X75Y125_SLICE_X115Y125_AO5),
.O6(CLBLL_R_X75Y125_SLICE_X115Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y125_SLICE_X115Y125_MUXF7A (
.I0(CLBLL_R_X75Y125_SLICE_X115Y125_BO6),
.I1(CLBLL_R_X75Y125_SLICE_X115Y125_AO6),
.O(CLBLL_R_X75Y125_SLICE_X115Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y126_SLICE_X114Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y126_SLICE_X114Y126_DO5),
.O6(CLBLL_R_X75Y126_SLICE_X114Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y126_SLICE_X114Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y126_SLICE_X114Y126_CO5),
.O6(CLBLL_R_X75Y126_SLICE_X114Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y126_SLICE_X114Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y126_SLICE_X114Y126_BO5),
.O6(CLBLL_R_X75Y126_SLICE_X114Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y126_SLICE_X114Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y126_SLICE_X114Y126_AO5),
.O6(CLBLL_R_X75Y126_SLICE_X114Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf8cbc83b380b08)
  ) CLBLL_R_X75Y126_SLICE_X115Y126_DLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.O5(CLBLL_R_X75Y126_SLICE_X115Y126_DO5),
.O6(CLBLL_R_X75Y126_SLICE_X115Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccaafff0ccaa00)
  ) CLBLL_R_X75Y126_SLICE_X115Y126_CLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I2(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.O5(CLBLL_R_X75Y126_SLICE_X115Y126_CO5),
.O6(CLBLL_R_X75Y126_SLICE_X115Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050dd88dd88)
  ) CLBLL_R_X75Y126_SLICE_X115Y126_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I2(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X75Y126_SLICE_X115Y126_BO5),
.O6(CLBLL_R_X75Y126_SLICE_X115Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLL_R_X75Y126_SLICE_X115Y126_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I2(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLL_R_X75Y126_SLICE_X115Y126_AO5),
.O6(CLBLL_R_X75Y126_SLICE_X115Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y126_SLICE_X115Y126_MUXF7A (
.I0(CLBLL_R_X75Y126_SLICE_X115Y126_BO6),
.I1(CLBLL_R_X75Y126_SLICE_X115Y126_AO6),
.O(CLBLL_R_X75Y126_SLICE_X115Y126_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y126_SLICE_X115Y126_MUXF7B (
.I0(CLBLL_R_X75Y126_SLICE_X115Y126_DO6),
.I1(CLBLL_R_X75Y126_SLICE_X115Y126_CO6),
.O(CLBLL_R_X75Y126_SLICE_X115Y126_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y127_SLICE_X114Y127_DO5),
.O6(CLBLL_R_X75Y127_SLICE_X114Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h56569a9a569a569a)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_CLUT (
.I0(CLBLM_L_X70Y122_SLICE_X104Y122_CO6),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(CLBLL_R_X75Y127_SLICE_X115Y127_F8MUX_O),
.I3(CLBLL_R_X75Y127_SLICE_X114Y127_F7AMUX_O),
.I4(CLBLM_L_X74Y127_SLICE_X113Y127_F7AMUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X75Y127_SLICE_X114Y127_CO5),
.O6(CLBLL_R_X75Y127_SLICE_X114Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_BLUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I1(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X75Y127_SLICE_X114Y127_BO5),
.O6(CLBLL_R_X75Y127_SLICE_X114Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0acfcffa0ac0c0)
  ) CLBLL_R_X75Y127_SLICE_X114Y127_ALUT (
.I0(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.O5(CLBLL_R_X75Y127_SLICE_X114Y127_AO5),
.O6(CLBLL_R_X75Y127_SLICE_X114Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y127_SLICE_X114Y127_MUXF7A (
.I0(CLBLL_R_X75Y127_SLICE_X114Y127_BO6),
.I1(CLBLL_R_X75Y127_SLICE_X114Y127_AO6),
.O(CLBLL_R_X75Y127_SLICE_X114Y127_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfa0afa0a)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_DLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X75Y127_SLICE_X115Y127_DO5),
.O6(CLBLL_R_X75Y127_SLICE_X115Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ffccaaf000ccaa)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_CLUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.O5(CLBLL_R_X75Y127_SLICE_X115Y127_CO5),
.O6(CLBLL_R_X75Y127_SLICE_X115Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf8ada85d580d08)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_BLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.O5(CLBLL_R_X75Y127_SLICE_X115Y127_BO5),
.O6(CLBLL_R_X75Y127_SLICE_X115Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLL_R_X75Y127_SLICE_X115Y127_ALUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I1(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLL_R_X75Y127_SLICE_X115Y127_AO5),
.O6(CLBLL_R_X75Y127_SLICE_X115Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y127_SLICE_X115Y127_MUXF7A (
.I0(CLBLL_R_X75Y127_SLICE_X115Y127_BO6),
.I1(CLBLL_R_X75Y127_SLICE_X115Y127_AO6),
.O(CLBLL_R_X75Y127_SLICE_X115Y127_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y127_SLICE_X115Y127_MUXF7B (
.I0(CLBLL_R_X75Y127_SLICE_X115Y127_DO6),
.I1(CLBLL_R_X75Y127_SLICE_X115Y127_CO6),
.O(CLBLL_R_X75Y127_SLICE_X115Y127_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X75Y127_SLICE_X115Y127_MUXF8 (
.I0(CLBLL_R_X75Y127_SLICE_X115Y127_F7BMUX_O),
.I1(CLBLL_R_X75Y127_SLICE_X115Y127_F7AMUX_O),
.O(CLBLL_R_X75Y127_SLICE_X115Y127_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbd97351eac86240)
  ) CLBLL_R_X75Y128_SLICE_X114Y128_DLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I5(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.O5(CLBLL_R_X75Y128_SLICE_X114Y128_DO5),
.O6(CLBLL_R_X75Y128_SLICE_X114Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ffaa5500)
  ) CLBLL_R_X75Y128_SLICE_X114Y128_CLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X75Y128_SLICE_X114Y128_CO5),
.O6(CLBLL_R_X75Y128_SLICE_X114Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe5eae0ef454a404)
  ) CLBLL_R_X75Y128_SLICE_X114Y128_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.O5(CLBLL_R_X75Y128_SLICE_X114Y128_BO5),
.O6(CLBLL_R_X75Y128_SLICE_X114Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffac0facf0ac00ac)
  ) CLBLL_R_X75Y128_SLICE_X114Y128_ALUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I1(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I5(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.O5(CLBLL_R_X75Y128_SLICE_X114Y128_AO5),
.O6(CLBLL_R_X75Y128_SLICE_X114Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y128_SLICE_X114Y128_MUXF7A (
.I0(CLBLL_R_X75Y128_SLICE_X114Y128_BO6),
.I1(CLBLL_R_X75Y128_SLICE_X114Y128_AO6),
.O(CLBLL_R_X75Y128_SLICE_X114Y128_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y128_SLICE_X114Y128_MUXF7B (
.I0(CLBLL_R_X75Y128_SLICE_X114Y128_DO6),
.I1(CLBLL_R_X75Y128_SLICE_X114Y128_CO6),
.O(CLBLL_R_X75Y128_SLICE_X114Y128_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X75Y128_SLICE_X114Y128_MUXF8 (
.I0(CLBLL_R_X75Y128_SLICE_X114Y128_F7BMUX_O),
.I1(CLBLL_R_X75Y128_SLICE_X114Y128_F7AMUX_O),
.O(CLBLL_R_X75Y128_SLICE_X114Y128_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X75Y128_SLICE_X115Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X75Y128_SLICE_X115Y128_DO5),
.O6(CLBLL_R_X75Y128_SLICE_X115Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fa55af02d2d7878)
  ) CLBLL_R_X75Y128_SLICE_X115Y128_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_F7AMUX_O),
.I2(CLBLL_L_X2Y123_SLICE_X0Y123_DO6),
.I3(CLBLL_R_X75Y128_SLICE_X115Y128_F7AMUX_O),
.I4(CLBLM_L_X76Y128_SLICE_X116Y128_F8MUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLL_R_X75Y128_SLICE_X115Y128_CO5),
.O6(CLBLL_R_X75Y128_SLICE_X115Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2ffe233e2cce200)
  ) CLBLL_R_X75Y128_SLICE_X115Y128_BLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I5(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.O5(CLBLL_R_X75Y128_SLICE_X115Y128_BO5),
.O6(CLBLL_R_X75Y128_SLICE_X115Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0aaffccf0aa00)
  ) CLBLL_R_X75Y128_SLICE_X115Y128_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I1(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.O5(CLBLL_R_X75Y128_SLICE_X115Y128_AO5),
.O6(CLBLL_R_X75Y128_SLICE_X115Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X75Y128_SLICE_X115Y128_MUXF7A (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_BO6),
.I1(CLBLL_R_X75Y128_SLICE_X115Y128_AO6),
.O(CLBLL_R_X75Y128_SLICE_X115Y128_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000be82be82)
  ) CLBLL_R_X77Y113_SLICE_X118Y113_DLUT (
.I0(LIOB33_X0Y151_IOB_X0Y152_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y113_SLICE_X118Y113_DO5),
.O6(CLBLL_R_X77Y113_SLICE_X118Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000caaccaac)
  ) CLBLL_R_X77Y113_SLICE_X118Y113_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_SING_X0Y150_IOB_X0Y150_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y113_SLICE_X118Y113_CO5),
.O6(CLBLL_R_X77Y113_SLICE_X118Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffed00edff480048)
  ) CLBLL_R_X77Y113_SLICE_X118Y113_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y151_IOB_X0Y151_I),
.O5(CLBLL_R_X77Y113_SLICE_X118Y113_BO5),
.O6(CLBLL_R_X77Y113_SLICE_X118Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f690f690)
  ) CLBLL_R_X77Y113_SLICE_X118Y113_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(LIOB33_X0Y155_IOB_X0Y156_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_SING_X105Y50_IOB_X1Y50_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y113_SLICE_X118Y113_AO5),
.O6(CLBLL_R_X77Y113_SLICE_X118Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X119Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X119Y113_DO5),
.O6(CLBLL_R_X77Y113_SLICE_X119Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X119Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X119Y113_CO5),
.O6(CLBLL_R_X77Y113_SLICE_X119Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X119Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X119Y113_BO5),
.O6(CLBLL_R_X77Y113_SLICE_X119Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y113_SLICE_X119Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y113_SLICE_X119Y113_AO5),
.O6(CLBLL_R_X77Y113_SLICE_X119Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y114_SLICE_X118Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y114_SLICE_X118Y114_DO5),
.O6(CLBLL_R_X77Y114_SLICE_X118Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y114_SLICE_X118Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y114_SLICE_X118Y114_CO5),
.O6(CLBLL_R_X77Y114_SLICE_X118Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000e4d8e4d8)
  ) CLBLL_R_X77Y114_SLICE_X118Y114_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_X0Y157_IOB_X0Y157_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(RIOB33_X105Y51_IOB_X1Y51_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y114_SLICE_X118Y114_BO5),
.O6(CLBLL_R_X77Y114_SLICE_X118Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc50ccf5cca0)
  ) CLBLL_R_X77Y114_SLICE_X118Y114_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y51_IOB_X1Y52_I),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(LIOB33_X0Y157_IOB_X0Y158_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLL_R_X77Y114_SLICE_X118Y114_AO5),
.O6(CLBLL_R_X77Y114_SLICE_X118Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y114_SLICE_X119Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y114_SLICE_X119Y114_DO5),
.O6(CLBLL_R_X77Y114_SLICE_X119Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y114_SLICE_X119Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y114_SLICE_X119Y114_CO5),
.O6(CLBLL_R_X77Y114_SLICE_X119Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y114_SLICE_X119Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y114_SLICE_X119Y114_BO5),
.O6(CLBLL_R_X77Y114_SLICE_X119Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y114_SLICE_X119Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y114_SLICE_X119Y114_AO5),
.O6(CLBLL_R_X77Y114_SLICE_X119Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y115_SLICE_X118Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y115_SLICE_X118Y115_DO5),
.O6(CLBLL_R_X77Y115_SLICE_X118Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y115_SLICE_X118Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y115_SLICE_X118Y115_CO5),
.O6(CLBLL_R_X77Y115_SLICE_X118Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y115_SLICE_X118Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y115_SLICE_X118Y115_BO5),
.O6(CLBLL_R_X77Y115_SLICE_X118Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f960f960)
  ) CLBLL_R_X77Y115_SLICE_X118Y115_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(LIOB33_X0Y159_IOB_X0Y159_I),
.I4(RIOB33_X105Y53_IOB_X1Y53_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y115_SLICE_X118Y115_AO5),
.O6(CLBLL_R_X77Y115_SLICE_X118Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y115_SLICE_X119Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y115_SLICE_X119Y115_DO5),
.O6(CLBLL_R_X77Y115_SLICE_X119Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y115_SLICE_X119Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y115_SLICE_X119Y115_CO5),
.O6(CLBLL_R_X77Y115_SLICE_X119Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y115_SLICE_X119Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y115_SLICE_X119Y115_BO5),
.O6(CLBLL_R_X77Y115_SLICE_X119Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y115_SLICE_X119Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y115_SLICE_X119Y115_AO5),
.O6(CLBLL_R_X77Y115_SLICE_X119Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbeebaa55144100)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_DLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y179_IOB_X0Y179_I),
.I4(RIOB33_X105Y189_IOB_X1Y189_I),
.I5(RIOB33_X105Y73_IOB_X1Y73_I),
.O5(CLBLL_R_X77Y122_SLICE_X118Y122_DO5),
.O6(CLBLL_R_X77Y122_SLICE_X118Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32ef23ce02ec20)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_CLUT (
.I0(RIOB33_X105Y195_IOB_X1Y196_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(RIOB33_X105Y95_IOB_X1Y96_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(LIOB33_X0Y201_IOB_X0Y202_I),
.O5(CLBLL_R_X77Y122_SLICE_X118Y122_CO5),
.O6(CLBLL_R_X77Y122_SLICE_X118Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffde3312edcc2100)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y177_IOB_X0Y178_I),
.I4(RIOB33_X105Y71_IOB_X1Y72_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_R_X77Y122_SLICE_X118Y122_BO5),
.O6(CLBLL_R_X77Y122_SLICE_X118Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc5acca5cc00)
  ) CLBLL_R_X77Y122_SLICE_X118Y122_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y89_IOB_X1Y89_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(LIOB33_X0Y195_IOB_X0Y195_I),
.I5(RIOB33_X105Y145_IOB_X1Y145_I),
.O5(CLBLL_R_X77Y122_SLICE_X118Y122_AO5),
.O6(CLBLL_R_X77Y122_SLICE_X118Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y122_SLICE_X119Y122_DO5),
.O6(CLBLL_R_X77Y122_SLICE_X119Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y122_SLICE_X119Y122_CO5),
.O6(CLBLL_R_X77Y122_SLICE_X119Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y122_SLICE_X119Y122_BO5),
.O6(CLBLL_R_X77Y122_SLICE_X119Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y122_SLICE_X119Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y122_SLICE_X119Y122_AO5),
.O6(CLBLL_R_X77Y122_SLICE_X119Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacfff00f00)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_DLUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I1(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X77Y125_SLICE_X118Y125_DO5),
.O6(CLBLL_R_X77Y125_SLICE_X118Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0aaaacccc)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_CLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X77Y125_SLICE_X118Y125_CO5),
.O6(CLBLL_R_X77Y125_SLICE_X118Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88fafa5050)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_BLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I2(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_R_X77Y125_SLICE_X118Y125_BO5),
.O6(CLBLL_R_X77Y125_SLICE_X118Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfadd5088fa8850)
  ) CLBLL_R_X77Y125_SLICE_X118Y125_ALUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.O5(CLBLL_R_X77Y125_SLICE_X118Y125_AO5),
.O6(CLBLL_R_X77Y125_SLICE_X118Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLL_R_X77Y125_SLICE_X118Y125_MUXF7A (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_BO6),
.I1(CLBLL_R_X77Y125_SLICE_X118Y125_AO6),
.O(CLBLL_R_X77Y125_SLICE_X118Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLL_R_X77Y125_SLICE_X118Y125_MUXF7B (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_DO6),
.I1(CLBLL_R_X77Y125_SLICE_X118Y125_CO6),
.O(CLBLL_R_X77Y125_SLICE_X118Y125_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLL_R_X77Y125_SLICE_X118Y125_MUXF8 (
.I0(CLBLL_R_X77Y125_SLICE_X118Y125_F7BMUX_O),
.I1(CLBLL_R_X77Y125_SLICE_X118Y125_F7AMUX_O),
.O(CLBLL_R_X77Y125_SLICE_X118Y125_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y125_SLICE_X119Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X119Y125_DO5),
.O6(CLBLL_R_X77Y125_SLICE_X119Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y125_SLICE_X119Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X119Y125_CO5),
.O6(CLBLL_R_X77Y125_SLICE_X119Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y125_SLICE_X119Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X119Y125_BO5),
.O6(CLBLL_R_X77Y125_SLICE_X119Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y125_SLICE_X119Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y125_SLICE_X119Y125_AO5),
.O6(CLBLL_R_X77Y125_SLICE_X119Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb800b8ffe200e2)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_DLUT (
.I0(LIOB33_SING_X0Y200_IOB_X0Y200_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(RIOB33_X105Y193_IOB_X1Y194_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(RIOB33_X105Y93_IOB_X1Y94_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLL_R_X77Y129_SLICE_X118Y129_DO5),
.O6(CLBLL_R_X77Y129_SLICE_X118Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffde00deff840084)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_CLUT (
.I0(LIOB33_X0Y85_IOB_X0Y85_I),
.I1(LIOB33_X0Y193_IOB_X0Y194_I),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(RIOB33_X105Y87_IOB_X1Y88_I),
.I5(RIOB33_X105Y143_IOB_X1Y144_I),
.O5(CLBLL_R_X77Y129_SLICE_X118Y129_CO5),
.O6(CLBLL_R_X77Y129_SLICE_X118Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d8e4d8e4)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_BLUT (
.I0(LIOB33_X0Y85_IOB_X0Y85_I),
.I1(LIOB33_X0Y201_IOB_X0Y201_I),
.I2(RIOB33_X105Y195_IOB_X1Y195_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(RIOB33_X105Y95_IOB_X1Y95_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y129_SLICE_X118Y129_BO5),
.O6(CLBLL_R_X77Y129_SLICE_X118Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0eebb2288)
  ) CLBLL_R_X77Y129_SLICE_X118Y129_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(RIOB33_X105Y69_IOB_X1Y69_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(LIOB33_X0Y175_IOB_X0Y175_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y129_SLICE_X118Y129_AO5),
.O6(CLBLL_R_X77Y129_SLICE_X118Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y129_SLICE_X119Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y129_SLICE_X119Y129_DO5),
.O6(CLBLL_R_X77Y129_SLICE_X119Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y129_SLICE_X119Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y129_SLICE_X119Y129_CO5),
.O6(CLBLL_R_X77Y129_SLICE_X119Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y129_SLICE_X119Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y129_SLICE_X119Y129_BO5),
.O6(CLBLL_R_X77Y129_SLICE_X119Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y129_SLICE_X119Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y129_SLICE_X119Y129_AO5),
.O6(CLBLL_R_X77Y129_SLICE_X119Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe200e2ffb800b8)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(LIOB33_X0Y177_IOB_X0Y177_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(RIOB33_X105Y71_IOB_X1Y71_I),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLL_R_X77Y130_SLICE_X118Y130_DO5),
.O6(CLBLL_R_X77Y130_SLICE_X118Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0bbf088f0eef022)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_CLUT (
.I0(LIOB33_X0Y203_IOB_X0Y203_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(RIOB33_X105Y97_IOB_X1Y97_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(RIOB33_X105Y197_IOB_X1Y197_I),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLL_R_X77Y130_SLICE_X118Y130_CO5),
.O6(CLBLL_R_X77Y130_SLICE_X118Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefbbaea54511040)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(RIOB33_X105Y187_IOB_X1Y188_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(LIOB33_X0Y169_IOB_X0Y169_I),
.I5(RIOB33_X105Y63_IOB_X1Y63_I),
.O5(CLBLL_R_X77Y130_SLICE_X118Y130_BO5),
.O6(CLBLL_R_X77Y130_SLICE_X118Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000be82be82)
  ) CLBLL_R_X77Y130_SLICE_X118Y130_ALUT (
.I0(LIOB33_X0Y183_IOB_X0Y183_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(RIOB33_X105Y193_IOB_X1Y193_I),
.I4(RIOB33_X105Y77_IOB_X1Y77_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y130_SLICE_X118Y130_AO5),
.O6(CLBLL_R_X77Y130_SLICE_X118Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y130_SLICE_X119Y130_DO5),
.O6(CLBLL_R_X77Y130_SLICE_X119Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y130_SLICE_X119Y130_CO5),
.O6(CLBLL_R_X77Y130_SLICE_X119Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y130_SLICE_X119Y130_BO5),
.O6(CLBLL_R_X77Y130_SLICE_X119Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y130_SLICE_X119Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y130_SLICE_X119Y130_AO5),
.O6(CLBLL_R_X77Y130_SLICE_X119Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaf0aaf0aacc)
  ) CLBLL_R_X77Y131_SLICE_X118Y131_DLUT (
.I0(RIOB33_X105Y69_IOB_X1Y70_I),
.I1(LIOB33_X0Y175_IOB_X0Y176_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(LIOB33_X0Y85_IOB_X0Y85_I),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLL_R_X77Y131_SLICE_X118Y131_DO5),
.O6(CLBLL_R_X77Y131_SLICE_X118Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000de84de84)
  ) CLBLL_R_X77Y131_SLICE_X118Y131_CLUT (
.I0(LIOB33_X0Y85_IOB_X0Y85_I),
.I1(LIOB33_X0Y195_IOB_X0Y196_I),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(RIOB33_X105Y89_IOB_X1Y90_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y131_SLICE_X118Y131_CO5),
.O6(CLBLL_R_X77Y131_SLICE_X118Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00d8d8e4e4)
  ) CLBLL_R_X77Y131_SLICE_X118Y131_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y189_IOB_X0Y189_I),
.I2(RIOB33_X105Y139_IOB_X1Y139_I),
.I3(RIOB33_X105Y83_IOB_X1Y83_I),
.I4(LIOB33_X0Y85_IOB_X0Y85_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y131_SLICE_X118Y131_BO5),
.O6(CLBLL_R_X77Y131_SLICE_X118Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccaaaacc)
  ) CLBLL_R_X77Y131_SLICE_X118Y131_ALUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(LIOB33_X0Y197_IOB_X0Y197_I),
.I2(RIOB33_X105Y91_IOB_X1Y91_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(LIOB33_X0Y85_IOB_X0Y85_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y131_SLICE_X118Y131_AO5),
.O6(CLBLL_R_X77Y131_SLICE_X118Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y131_SLICE_X119Y131_DO5),
.O6(CLBLL_R_X77Y131_SLICE_X119Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y131_SLICE_X119Y131_CO5),
.O6(CLBLL_R_X77Y131_SLICE_X119Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y131_SLICE_X119Y131_BO5),
.O6(CLBLL_R_X77Y131_SLICE_X119Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y131_SLICE_X119Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y131_SLICE_X119Y131_AO5),
.O6(CLBLL_R_X77Y131_SLICE_X119Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y133_SLICE_X118Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y133_SLICE_X118Y133_DO5),
.O6(CLBLL_R_X77Y133_SLICE_X118Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y133_SLICE_X118Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y133_SLICE_X118Y133_CO5),
.O6(CLBLL_R_X77Y133_SLICE_X118Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000be82be82)
  ) CLBLL_R_X77Y133_SLICE_X118Y133_BLUT (
.I0(LIOB33_X0Y181_IOB_X0Y182_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(RIOB33_X105Y191_IOB_X1Y192_I),
.I4(RIOB33_X105Y75_IOB_X1Y76_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y133_SLICE_X118Y133_BO5),
.O6(CLBLL_R_X77Y133_SLICE_X118Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ed48ed48)
  ) CLBLL_R_X77Y133_SLICE_X118Y133_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y141_IOB_X1Y141_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y191_IOB_X0Y191_I),
.I4(RIOB33_X105Y85_IOB_X1Y85_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLL_R_X77Y133_SLICE_X118Y133_AO5),
.O6(CLBLL_R_X77Y133_SLICE_X118Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y133_SLICE_X119Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y133_SLICE_X119Y133_DO5),
.O6(CLBLL_R_X77Y133_SLICE_X119Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y133_SLICE_X119Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y133_SLICE_X119Y133_CO5),
.O6(CLBLL_R_X77Y133_SLICE_X119Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y133_SLICE_X119Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y133_SLICE_X119Y133_BO5),
.O6(CLBLL_R_X77Y133_SLICE_X119Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X77Y133_SLICE_X119Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X77Y133_SLICE_X119Y133_AO5),
.O6(CLBLL_R_X77Y133_SLICE_X119Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y123_SLICE_X122Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y123_SLICE_X122Y123_DO5),
.O6(CLBLL_R_X79Y123_SLICE_X122Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y123_SLICE_X122Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y123_SLICE_X122Y123_CO5),
.O6(CLBLL_R_X79Y123_SLICE_X122Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0dd88f0f0ee44)
  ) CLBLL_R_X79Y123_SLICE_X122Y123_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y185_IOB_X0Y186_I),
.I2(RIOB33_X105Y79_IOB_X1Y80_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(LIOB33_X0Y83_IOB_X0Y83_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLL_R_X79Y123_SLICE_X122Y123_BO5),
.O6(CLBLL_R_X79Y123_SLICE_X122Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc5cac0cfcac5c0)
  ) CLBLL_R_X79Y123_SLICE_X122Y123_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y61_IOB_X1Y61_I),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(LIOB33_X0Y167_IOB_X0Y167_I),
.I4(RIOB33_X105Y123_IOB_X1Y123_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLL_R_X79Y123_SLICE_X122Y123_AO5),
.O6(CLBLL_R_X79Y123_SLICE_X122Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y123_SLICE_X123Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y123_SLICE_X123Y123_DO5),
.O6(CLBLL_R_X79Y123_SLICE_X123Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y123_SLICE_X123Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y123_SLICE_X123Y123_CO5),
.O6(CLBLL_R_X79Y123_SLICE_X123Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y123_SLICE_X123Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y123_SLICE_X123Y123_BO5),
.O6(CLBLL_R_X79Y123_SLICE_X123Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y123_SLICE_X123Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y123_SLICE_X123Y123_AO5),
.O6(CLBLL_R_X79Y123_SLICE_X123Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y124_SLICE_X122Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y124_SLICE_X122Y124_DO5),
.O6(CLBLL_R_X79Y124_SLICE_X122Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcacacfc0cacac0)
  ) CLBLL_R_X79Y124_SLICE_X122Y124_CLUT (
.I0(RIOB33_X105Y127_IOB_X1Y127_I),
.I1(RIOB33_X105Y65_IOB_X1Y66_I),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(LIOB33_X0Y171_IOB_X0Y172_I),
.O5(CLBLL_R_X79Y124_SLICE_X122Y124_CO5),
.O6(CLBLL_R_X79Y124_SLICE_X122Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0ef404fd0df808)
  ) CLBLL_R_X79Y124_SLICE_X122Y124_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(RIOB33_X105Y67_IOB_X1Y67_I),
.I4(LIOB33_X0Y173_IOB_X0Y173_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLL_R_X79Y124_SLICE_X122Y124_BO5),
.O6(CLBLL_R_X79Y124_SLICE_X122Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc5cac0cfcac5c0)
  ) CLBLL_R_X79Y124_SLICE_X122Y124_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y61_IOB_X1Y62_I),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(LIOB33_X0Y167_IOB_X0Y168_I),
.I4(RIOB33_X105Y123_IOB_X1Y124_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLL_R_X79Y124_SLICE_X122Y124_AO5),
.O6(CLBLL_R_X79Y124_SLICE_X122Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y124_SLICE_X123Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y124_SLICE_X123Y124_DO5),
.O6(CLBLL_R_X79Y124_SLICE_X123Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y124_SLICE_X123Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y124_SLICE_X123Y124_CO5),
.O6(CLBLL_R_X79Y124_SLICE_X123Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y124_SLICE_X123Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y124_SLICE_X123Y124_BO5),
.O6(CLBLL_R_X79Y124_SLICE_X123Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y124_SLICE_X123Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y124_SLICE_X123Y124_AO5),
.O6(CLBLL_R_X79Y124_SLICE_X123Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y125_SLICE_X122Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y125_SLICE_X122Y125_DO5),
.O6(CLBLL_R_X79Y125_SLICE_X122Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y125_SLICE_X122Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y125_SLICE_X122Y125_CO5),
.O6(CLBLL_R_X79Y125_SLICE_X122Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y125_SLICE_X122Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y125_SLICE_X122Y125_BO5),
.O6(CLBLL_R_X79Y125_SLICE_X122Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31ec20fe32dc10)
  ) CLBLL_R_X79Y125_SLICE_X122Y125_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(LIOB33_X0Y169_IOB_X0Y170_I),
.I3(RIOB33_X105Y63_IOB_X1Y64_I),
.I4(RIOB33_X105Y125_IOB_X1Y125_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLL_R_X79Y125_SLICE_X122Y125_AO5),
.O6(CLBLL_R_X79Y125_SLICE_X122Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y125_SLICE_X123Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y125_SLICE_X123Y125_DO5),
.O6(CLBLL_R_X79Y125_SLICE_X123Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y125_SLICE_X123Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y125_SLICE_X123Y125_CO5),
.O6(CLBLL_R_X79Y125_SLICE_X123Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y125_SLICE_X123Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y125_SLICE_X123Y125_BO5),
.O6(CLBLL_R_X79Y125_SLICE_X123Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_R_X79Y125_SLICE_X123Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_R_X79Y125_SLICE_X123Y125_AO5),
.O6(CLBLL_R_X79Y125_SLICE_X123Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y118_SLICE_X66Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y118_SLICE_X66Y118_DO5),
.O6(CLBLM_L_X44Y118_SLICE_X66Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y118_SLICE_X66Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y118_SLICE_X66Y118_CO5),
.O6(CLBLM_L_X44Y118_SLICE_X66Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y118_SLICE_X66Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y118_SLICE_X66Y118_BO5),
.O6(CLBLM_L_X44Y118_SLICE_X66Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fff0ff00fff0)
  ) CLBLM_L_X44Y118_SLICE_X66Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(LIOB33_X0Y79_IOB_X0Y80_I),
.I5(1'b1),
.O5(CLBLM_L_X44Y118_SLICE_X66Y118_AO5),
.O6(CLBLM_L_X44Y118_SLICE_X66Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y118_SLICE_X67Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y118_SLICE_X67Y118_DO5),
.O6(CLBLM_L_X44Y118_SLICE_X67Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y118_SLICE_X67Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y118_SLICE_X67Y118_CO5),
.O6(CLBLM_L_X44Y118_SLICE_X67Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y118_SLICE_X67Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y118_SLICE_X67Y118_BO5),
.O6(CLBLM_L_X44Y118_SLICE_X67Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X44Y118_SLICE_X67Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X44Y118_SLICE_X67Y118_AO5),
.O6(CLBLM_L_X44Y118_SLICE_X67Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y116_SLICE_X70Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y116_SLICE_X70Y116_DO5),
.O6(CLBLM_L_X46Y116_SLICE_X70Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y116_SLICE_X70Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y116_SLICE_X70Y116_CO5),
.O6(CLBLM_L_X46Y116_SLICE_X70Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_L_X46Y116_SLICE_X70Y116_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLM_L_X46Y116_SLICE_X70Y116_BO5),
.O6(CLBLM_L_X46Y116_SLICE_X70Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_L_X46Y116_SLICE_X70Y116_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLM_L_X46Y116_SLICE_X70Y116_AO5),
.O6(CLBLM_L_X46Y116_SLICE_X70Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y116_SLICE_X71Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y116_SLICE_X71Y116_DO5),
.O6(CLBLM_L_X46Y116_SLICE_X71Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y116_SLICE_X71Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y116_SLICE_X71Y116_CO5),
.O6(CLBLM_L_X46Y116_SLICE_X71Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y116_SLICE_X71Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y116_SLICE_X71Y116_BO5),
.O6(CLBLM_L_X46Y116_SLICE_X71Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X46Y116_SLICE_X71Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X46Y116_SLICE_X71Y116_AO5),
.O6(CLBLM_L_X46Y116_SLICE_X71Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y116_SLICE_X84Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X56Y116_SLICE_X84Y116_CO6),
.Q(CLBLM_L_X56Y116_SLICE_X84Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X56Y116_SLICE_X84Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X56Y116_SLICE_X84Y116_AO6),
.Q(CLBLM_L_X56Y116_SLICE_X84Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y116_SLICE_X84Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y116_SLICE_X84Y116_DO5),
.O6(CLBLM_L_X56Y116_SLICE_X84Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000cccaccca)
  ) CLBLM_L_X56Y116_SLICE_X84Y116_CLUT (
.I0(CLBLM_L_X56Y116_SLICE_X84Y116_BQ),
.I1(CLBLM_L_X56Y116_SLICE_X84Y116_AQ),
.I2(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I4(RIOB33_X105Y165_IOB_X1Y165_I),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLM_L_X56Y116_SLICE_X84Y116_CO5),
.O6(CLBLM_L_X56Y116_SLICE_X84Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e4f0ddf0e4f088)
  ) CLBLM_L_X56Y116_SLICE_X84Y116_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLM_L_X56Y116_SLICE_X84Y116_BQ),
.I2(CLBLM_L_X56Y116_SLICE_X84Y116_AQ),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(LIOB33_X0Y55_IOB_X0Y55_I),
.O5(CLBLM_L_X56Y116_SLICE_X84Y116_BO5),
.O6(CLBLM_L_X56Y116_SLICE_X84Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e1ff0f0f1e0)
  ) CLBLM_L_X56Y116_SLICE_X84Y116_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(CLBLM_L_X56Y116_SLICE_X84Y116_AQ),
.I3(CLBLM_L_X56Y116_SLICE_X84Y116_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_R_X71Y116_SLICE_X107Y116_BO6),
.O5(CLBLM_L_X56Y116_SLICE_X84Y116_AO5),
.O6(CLBLM_L_X56Y116_SLICE_X84Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y116_SLICE_X85Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y116_SLICE_X85Y116_DO5),
.O6(CLBLM_L_X56Y116_SLICE_X85Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y116_SLICE_X85Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y116_SLICE_X85Y116_CO5),
.O6(CLBLM_L_X56Y116_SLICE_X85Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y116_SLICE_X85Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y116_SLICE_X85Y116_BO5),
.O6(CLBLM_L_X56Y116_SLICE_X85Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X56Y116_SLICE_X85Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X56Y116_SLICE_X85Y116_AO5),
.O6(CLBLM_L_X56Y116_SLICE_X85Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y119_SLICE_X102Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y119_SLICE_X102Y119_DO5),
.O6(CLBLM_L_X68Y119_SLICE_X102Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y119_SLICE_X102Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y119_SLICE_X102Y119_CO5),
.O6(CLBLM_L_X68Y119_SLICE_X102Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y119_SLICE_X102Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y119_SLICE_X102Y119_BO5),
.O6(CLBLM_L_X68Y119_SLICE_X102Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y119_SLICE_X102Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y119_SLICE_X102Y119_AO5),
.O6(CLBLM_L_X68Y119_SLICE_X102Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X68Y119_SLICE_X103Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X68Y119_SLICE_X103Y119_DO5),
.O6(CLBLM_L_X68Y119_SLICE_X103Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h994e69a54b9c26da)
  ) CLBLM_L_X68Y119_SLICE_X103Y119_CLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_CO6),
.I1(CLBLM_L_X70Y117_SLICE_X105Y117_AO6),
.I2(CLBLL_R_X73Y121_SLICE_X110Y121_CO6),
.I3(CLBLM_L_X72Y114_SLICE_X109Y114_CO6),
.I4(CLBLM_L_X72Y118_SLICE_X108Y118_DO6),
.I5(CLBLM_L_X72Y118_SLICE_X108Y118_CO6),
.O5(CLBLM_L_X68Y119_SLICE_X103Y119_CO5),
.O6(CLBLM_L_X68Y119_SLICE_X103Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6dc3c1799a699a26)
  ) CLBLM_L_X68Y119_SLICE_X103Y119_BLUT (
.I0(CLBLM_L_X72Y114_SLICE_X109Y114_CO6),
.I1(CLBLL_R_X73Y121_SLICE_X110Y121_CO6),
.I2(CLBLM_L_X72Y118_SLICE_X108Y118_DO6),
.I3(CLBLM_L_X72Y118_SLICE_X108Y118_CO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_CO6),
.I5(CLBLM_L_X70Y117_SLICE_X105Y117_AO6),
.O5(CLBLM_L_X68Y119_SLICE_X103Y119_BO5),
.O6(CLBLM_L_X68Y119_SLICE_X103Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h61971ed23e61e11e)
  ) CLBLM_L_X68Y119_SLICE_X103Y119_ALUT (
.I0(CLBLM_L_X72Y114_SLICE_X109Y114_CO6),
.I1(CLBLL_R_X73Y121_SLICE_X110Y121_CO6),
.I2(CLBLM_L_X72Y118_SLICE_X108Y118_DO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_CO6),
.I4(CLBLM_L_X72Y118_SLICE_X108Y118_CO6),
.I5(CLBLM_L_X70Y117_SLICE_X105Y117_AO6),
.O5(CLBLM_L_X68Y119_SLICE_X103Y119_AO5),
.O6(CLBLM_L_X68Y119_SLICE_X103Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y117_SLICE_X104Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y117_SLICE_X104Y117_DO5),
.O6(CLBLM_L_X70Y117_SLICE_X104Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y117_SLICE_X104Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y117_SLICE_X104Y117_CO5),
.O6(CLBLM_L_X70Y117_SLICE_X104Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y117_SLICE_X104Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y117_SLICE_X104Y117_BO5),
.O6(CLBLM_L_X70Y117_SLICE_X104Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y117_SLICE_X104Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y117_SLICE_X104Y117_AO5),
.O6(CLBLM_L_X70Y117_SLICE_X104Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y117_SLICE_X105Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y117_SLICE_X105Y117_DO5),
.O6(CLBLM_L_X70Y117_SLICE_X105Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y117_SLICE_X105Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y117_SLICE_X105Y117_CO5),
.O6(CLBLM_L_X70Y117_SLICE_X105Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y117_SLICE_X105Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y117_SLICE_X105Y117_BO5),
.O6(CLBLM_L_X70Y117_SLICE_X105Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fa52d2d5af07878)
  ) CLBLM_L_X70Y117_SLICE_X105Y117_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLL_R_X71Y117_SLICE_X106Y117_F7AMUX_O),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I3(CLBLL_R_X71Y117_SLICE_X106Y117_F7BMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_R_X71Y116_SLICE_X106Y116_F8MUX_O),
.O5(CLBLM_L_X70Y117_SLICE_X105Y117_AO5),
.O6(CLBLM_L_X70Y117_SLICE_X105Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y119_SLICE_X104Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y119_SLICE_X104Y119_AO6),
.Q(CLBLM_L_X70Y119_SLICE_X104Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y119_SLICE_X104Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X104Y119_DO5),
.O6(CLBLM_L_X70Y119_SLICE_X104Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbc41ca3d623d7e81)
  ) CLBLM_L_X70Y119_SLICE_X104Y119_CLUT (
.I0(CLBLM_L_X70Y117_SLICE_X105Y117_AO6),
.I1(CLBLM_L_X72Y114_SLICE_X109Y114_CO6),
.I2(CLBLM_L_X72Y118_SLICE_X108Y118_DO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_CO6),
.I4(CLBLL_R_X73Y121_SLICE_X110Y121_CO6),
.I5(CLBLM_L_X72Y118_SLICE_X108Y118_CO6),
.O5(CLBLM_L_X70Y119_SLICE_X104Y119_CO5),
.O6(CLBLM_L_X70Y119_SLICE_X104Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccd8ccf5ccd8cca0)
  ) CLBLM_L_X70Y119_SLICE_X104Y119_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLL_R_X71Y119_SLICE_X106Y119_AQ),
.I2(CLBLM_L_X70Y119_SLICE_X104Y119_AQ),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(RIOB33_SING_X105Y150_IOB_X1Y150_I),
.O5(CLBLM_L_X70Y119_SLICE_X104Y119_BO5),
.O6(CLBLM_L_X70Y119_SLICE_X104Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff01fdff00fe02)
  ) CLBLM_L_X70Y119_SLICE_X104Y119_ALUT (
.I0(CLBLM_L_X70Y119_SLICE_X104Y119_BO6),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(CLBLL_R_X71Y119_SLICE_X106Y119_AQ),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_R_X71Y119_SLICE_X106Y119_CO6),
.O5(CLBLM_L_X70Y119_SLICE_X104Y119_AO5),
.O6(CLBLM_L_X70Y119_SLICE_X104Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y119_SLICE_X105Y119_CO6),
.Q(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y119_SLICE_X105Y119_AO6),
.Q(CLBLM_L_X70Y119_SLICE_X105Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y119_SLICE_X105Y119_DO5),
.O6(CLBLM_L_X70Y119_SLICE_X105Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafeba55005410)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_CLUT (
.I0(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I2(CLBLM_L_X70Y119_SLICE_X105Y119_BQ),
.I3(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.I4(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I5(RIOB33_X105Y177_IOB_X1Y177_I),
.O5(CLBLM_L_X70Y119_SLICE_X105Y119_CO5),
.O6(CLBLM_L_X70Y119_SLICE_X105Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffedffe8004d0048)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLM_L_X70Y119_SLICE_X105Y119_BQ),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(RIOB33_X105Y175_IOB_X1Y176_I),
.I5(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.O5(CLBLM_L_X70Y119_SLICE_X105Y119_BO5),
.O6(CLBLM_L_X70Y119_SLICE_X105Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555457aaaaaba8)
  ) CLBLM_L_X70Y119_SLICE_X105Y119_ALUT (
.I0(CLBLM_L_X70Y119_SLICE_X105Y119_AQ),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(CLBLM_L_X70Y119_SLICE_X105Y119_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLL_R_X71Y116_SLICE_X107Y116_CO6),
.O5(CLBLM_L_X70Y119_SLICE_X105Y119_AO5),
.O6(CLBLM_L_X70Y119_SLICE_X105Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y121_SLICE_X104Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y123_SLICE_X104Y123_BO6),
.Q(CLBLM_L_X70Y121_SLICE_X104Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y121_SLICE_X104Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y121_SLICE_X104Y121_DO6),
.Q(CLBLM_L_X70Y121_SLICE_X104Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y121_SLICE_X104Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y121_SLICE_X104Y121_BO6),
.Q(CLBLM_L_X70Y121_SLICE_X104Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y121_SLICE_X104Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y121_SLICE_X104Y121_AO6),
.Q(CLBLM_L_X70Y121_SLICE_X104Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaff00acac)
  ) CLBLM_L_X70Y121_SLICE_X104Y121_DLUT (
.I0(CLBLM_L_X70Y121_SLICE_X104Y121_BQ),
.I1(CLBLM_L_X70Y121_SLICE_X104Y121_CQ),
.I2(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I3(RIOB33_X105Y179_IOB_X1Y179_I),
.I4(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.O5(CLBLM_L_X70Y121_SLICE_X104Y121_DO5),
.O6(CLBLM_L_X70Y121_SLICE_X104Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaccfacc0)
  ) CLBLM_L_X70Y121_SLICE_X104Y121_CLUT (
.I0(CLBLM_L_X70Y121_SLICE_X104Y121_BQ),
.I1(CLBLM_L_X70Y121_SLICE_X104Y121_CQ),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(RIOB33_X105Y177_IOB_X1Y178_I),
.I5(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.O5(CLBLM_L_X70Y121_SLICE_X104Y121_CO5),
.O6(CLBLM_L_X70Y121_SLICE_X104Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33323337cccdccc8)
  ) CLBLM_L_X70Y121_SLICE_X104Y121_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(CLBLM_L_X70Y121_SLICE_X104Y121_BQ),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(CLBLM_L_X70Y121_SLICE_X104Y121_CO6),
.I5(CLBLM_L_X72Y120_SLICE_X108Y120_CO6),
.O5(CLBLM_L_X70Y121_SLICE_X104Y121_BO5),
.O6(CLBLM_L_X70Y121_SLICE_X104Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f1bf0f0f0e4)
  ) CLBLM_L_X70Y121_SLICE_X104Y121_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(CLBLM_L_X70Y123_SLICE_X104Y123_AO6),
.I2(CLBLM_L_X70Y121_SLICE_X104Y121_AQ),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLL_R_X71Y119_SLICE_X106Y119_BO6),
.O5(CLBLM_L_X70Y121_SLICE_X104Y121_AO5),
.O6(CLBLM_L_X70Y121_SLICE_X104Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y121_SLICE_X105Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y121_SLICE_X105Y121_CO6),
.Q(CLBLM_L_X70Y121_SLICE_X105Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y121_SLICE_X105Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y121_SLICE_X105Y121_AO6),
.Q(CLBLM_L_X70Y121_SLICE_X105Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y121_SLICE_X105Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y121_SLICE_X105Y121_DO5),
.O6(CLBLM_L_X70Y121_SLICE_X105Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfffa000a)
  ) CLBLM_L_X70Y121_SLICE_X105Y121_CLUT (
.I0(CLBLM_L_X70Y121_SLICE_X105Y121_BQ),
.I1(RIOB33_X105Y175_IOB_X1Y175_I),
.I2(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I4(CLBLM_L_X70Y121_SLICE_X105Y121_AQ),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLM_L_X70Y121_SLICE_X105Y121_CO5),
.O6(CLBLM_L_X70Y121_SLICE_X105Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffedffe8004d0048)
  ) CLBLM_L_X70Y121_SLICE_X105Y121_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLM_L_X70Y121_SLICE_X105Y121_BQ),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(RIOB33_X105Y173_IOB_X1Y174_I),
.I5(CLBLM_L_X70Y121_SLICE_X105Y121_AQ),
.O5(CLBLM_L_X70Y121_SLICE_X105Y121_BO5),
.O6(CLBLM_L_X70Y121_SLICE_X105Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f1df0f0f0e2)
  ) CLBLM_L_X70Y121_SLICE_X105Y121_ALUT (
.I0(CLBLM_L_X70Y121_SLICE_X105Y121_BO6),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLM_L_X70Y121_SLICE_X105Y121_AQ),
.I3(LIOB33_X0Y79_IOB_X0Y80_I),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLL_R_X71Y116_SLICE_X107Y116_DO6),
.O5(CLBLM_L_X70Y121_SLICE_X105Y121_AO5),
.O6(CLBLM_L_X70Y121_SLICE_X105Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y122_SLICE_X104Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y122_SLICE_X104Y122_CO6),
.Q(CLBLM_L_X70Y122_SLICE_X104Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y122_SLICE_X104Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y122_SLICE_X104Y122_AO6),
.Q(CLBLM_L_X70Y122_SLICE_X104Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y122_SLICE_X104Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y122_SLICE_X104Y122_DO5),
.O6(CLBLM_L_X70Y122_SLICE_X104Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfcfa0c0a)
  ) CLBLM_L_X70Y122_SLICE_X104Y122_CLUT (
.I0(CLBLM_L_X70Y122_SLICE_X104Y122_BQ),
.I1(CLBLM_L_X70Y122_SLICE_X104Y122_AQ),
.I2(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I4(RIOB33_X105Y173_IOB_X1Y173_I),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.O5(CLBLM_L_X70Y122_SLICE_X104Y122_CO5),
.O6(CLBLM_L_X70Y122_SLICE_X104Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e4e4e4e4f5a0)
  ) CLBLM_L_X70Y122_SLICE_X104Y122_BLUT (
.I0(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I1(CLBLM_L_X70Y122_SLICE_X104Y122_BQ),
.I2(CLBLM_L_X70Y122_SLICE_X104Y122_AQ),
.I3(RIOB33_X105Y171_IOB_X1Y172_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLM_L_X70Y122_SLICE_X104Y122_BO5),
.O6(CLBLM_L_X70Y122_SLICE_X104Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e1ff0f0f1e0)
  ) CLBLM_L_X70Y122_SLICE_X104Y122_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(CLBLM_L_X70Y122_SLICE_X104Y122_AQ),
.I3(CLBLM_L_X70Y122_SLICE_X104Y122_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLM_L_X70Y119_SLICE_X104Y119_CO6),
.O5(CLBLM_L_X70Y122_SLICE_X104Y122_AO5),
.O6(CLBLM_L_X70Y122_SLICE_X104Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y122_SLICE_X105Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y122_SLICE_X105Y122_DO5),
.O6(CLBLM_L_X70Y122_SLICE_X105Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y122_SLICE_X105Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y122_SLICE_X105Y122_CO5),
.O6(CLBLM_L_X70Y122_SLICE_X105Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y122_SLICE_X105Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y122_SLICE_X105Y122_BO5),
.O6(CLBLM_L_X70Y122_SLICE_X105Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y122_SLICE_X105Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y122_SLICE_X105Y122_AO5),
.O6(CLBLM_L_X70Y122_SLICE_X105Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y123_SLICE_X104Y123_DO5),
.O6(CLBLM_L_X70Y123_SLICE_X104Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y123_SLICE_X104Y123_CO5),
.O6(CLBLM_L_X70Y123_SLICE_X104Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfffa000a)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_BLUT (
.I0(CLBLM_L_X70Y121_SLICE_X104Y121_DQ),
.I1(RIOB33_X105Y167_IOB_X1Y167_I),
.I2(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(CLBLM_L_X70Y121_SLICE_X104Y121_AQ),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLM_L_X70Y123_SLICE_X104Y123_BO5),
.O6(CLBLM_L_X70Y123_SLICE_X104Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa000affac00ac)
  ) CLBLM_L_X70Y123_SLICE_X104Y123_ALUT (
.I0(CLBLM_L_X70Y121_SLICE_X104Y121_DQ),
.I1(RIOB33_X105Y165_IOB_X1Y166_I),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(CLBLM_L_X70Y121_SLICE_X104Y121_AQ),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLM_L_X70Y123_SLICE_X104Y123_AO5),
.O6(CLBLM_L_X70Y123_SLICE_X104Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y123_SLICE_X105Y123_CO6),
.Q(CLBLM_L_X70Y123_SLICE_X105Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y123_SLICE_X105Y123_AO6),
.Q(CLBLM_L_X70Y123_SLICE_X105Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y123_SLICE_X105Y123_DO6),
.Q(CLBLM_L_X70Y123_SLICE_X105Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c5a)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_DLUT (
.I0(CLBLM_L_X70Y124_SLICE_X105Y124_AO6),
.I1(CLBLM_L_X70Y124_SLICE_X105Y124_AQ),
.I2(CLBLL_R_X71Y120_SLICE_X107Y120_DO6),
.I3(LIOB33_X0Y81_IOB_X0Y82_I),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(LIOB33_X0Y79_IOB_X0Y80_I),
.O5(CLBLM_L_X70Y123_SLICE_X105Y123_DO5),
.O6(CLBLM_L_X70Y123_SLICE_X105Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeccdc33320010)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_CLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I1(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I2(CLBLM_L_X70Y123_SLICE_X105Y123_BQ),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(CLBLM_L_X70Y123_SLICE_X105Y123_AQ),
.I5(RIOB33_X105Y169_IOB_X1Y169_I),
.O5(CLBLM_L_X70Y123_SLICE_X105Y123_CO5),
.O6(CLBLM_L_X70Y123_SLICE_X105Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaacaaacaacfaac0)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_BLUT (
.I0(CLBLM_L_X70Y123_SLICE_X105Y123_AQ),
.I1(CLBLM_L_X70Y123_SLICE_X105Y123_BQ),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(RIOB33_X105Y167_IOB_X1Y168_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLM_L_X70Y123_SLICE_X105Y123_BO5),
.O6(CLBLM_L_X70Y123_SLICE_X105Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa5457aba8)
  ) CLBLM_L_X70Y123_SLICE_X105Y123_ALUT (
.I0(CLBLM_L_X70Y123_SLICE_X105Y123_AQ),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(CLBLM_L_X70Y123_SLICE_X105Y123_BO6),
.I4(CLBLL_R_X73Y122_SLICE_X110Y122_CO6),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLM_L_X70Y123_SLICE_X105Y123_AO5),
.O6(CLBLM_L_X70Y123_SLICE_X105Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y124_SLICE_X104Y124_CO6),
.Q(CLBLM_L_X70Y124_SLICE_X104Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y124_SLICE_X104Y124_AO6),
.Q(CLBLM_L_X70Y124_SLICE_X104Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y124_SLICE_X104Y124_DO5),
.O6(CLBLM_L_X70Y124_SLICE_X104Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfdfcf80c0d0c08)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_CLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I1(CLBLM_L_X70Y124_SLICE_X104Y124_AQ),
.I2(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(CLBLM_L_X70Y124_SLICE_X104Y124_BQ),
.I5(RIOB33_X105Y161_IOB_X1Y161_I),
.O5(CLBLM_L_X70Y124_SLICE_X104Y124_CO5),
.O6(CLBLM_L_X70Y124_SLICE_X104Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffca000c00ca)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_BLUT (
.I0(RIOB33_X105Y159_IOB_X1Y160_I),
.I1(CLBLM_L_X70Y124_SLICE_X104Y124_BQ),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(CLBLM_L_X70Y124_SLICE_X104Y124_AQ),
.O5(CLBLM_L_X70Y124_SLICE_X104Y124_BO5),
.O6(CLBLM_L_X70Y124_SLICE_X104Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00e1ff1e0)
  ) CLBLM_L_X70Y124_SLICE_X104Y124_ALUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(LIOB33_X0Y79_IOB_X0Y80_I),
.I2(CLBLM_L_X70Y124_SLICE_X104Y124_AQ),
.I3(CLBLM_L_X70Y124_SLICE_X104Y124_BO6),
.I4(CLBLL_R_X73Y122_SLICE_X110Y122_AO6),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLM_L_X70Y124_SLICE_X104Y124_AO5),
.O6(CLBLM_L_X70Y124_SLICE_X104Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y124_SLICE_X105Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.Q(CLBLM_L_X70Y124_SLICE_X105Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y124_SLICE_X105Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y124_SLICE_X105Y124_DO5),
.O6(CLBLM_L_X70Y124_SLICE_X105Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y124_SLICE_X105Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y124_SLICE_X105Y124_CO5),
.O6(CLBLM_L_X70Y124_SLICE_X105Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8bbb8b8b888)
  ) CLBLM_L_X70Y124_SLICE_X105Y124_BLUT (
.I0(RIOB33_X105Y183_IOB_X1Y183_I),
.I1(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I2(CLBLM_L_X70Y124_SLICE_X105Y124_AQ),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I5(CLBLM_L_X70Y123_SLICE_X105Y123_CQ),
.O5(CLBLM_L_X70Y124_SLICE_X105Y124_BO5),
.O6(CLBLM_L_X70Y124_SLICE_X105Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f3e2f0c0c0e2)
  ) CLBLM_L_X70Y124_SLICE_X105Y124_ALUT (
.I0(RIOB33_X105Y181_IOB_X1Y182_I),
.I1(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I2(CLBLM_L_X70Y124_SLICE_X105Y124_AQ),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(CLBLM_L_X70Y123_SLICE_X105Y123_CQ),
.O5(CLBLM_L_X70Y124_SLICE_X105Y124_AO5),
.O6(CLBLM_L_X70Y124_SLICE_X105Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y127_SLICE_X104Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y127_SLICE_X104Y127_DO6),
.Q(CLBLM_L_X70Y127_SLICE_X104Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y127_SLICE_X104Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y127_SLICE_X104Y127_AO6),
.Q(CLBLM_L_X70Y127_SLICE_X104Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y127_SLICE_X104Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y127_SLICE_X104Y127_BO6),
.Q(CLBLM_L_X70Y127_SLICE_X104Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0f0cc)
  ) CLBLM_L_X70Y127_SLICE_X104Y127_DLUT (
.I0(RIOB33_X105Y185_IOB_X1Y185_I),
.I1(CLBLM_L_X70Y127_SLICE_X104Y127_CQ),
.I2(CLBLM_L_X70Y127_SLICE_X104Y127_AQ),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I4(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLM_L_X70Y127_SLICE_X104Y127_DO5),
.O6(CLBLM_L_X70Y127_SLICE_X104Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0e4e4f0f0dd88)
  ) CLBLM_L_X70Y127_SLICE_X104Y127_CLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLM_L_X70Y127_SLICE_X104Y127_CQ),
.I2(CLBLM_L_X70Y127_SLICE_X104Y127_AQ),
.I3(RIOB33_X105Y183_IOB_X1Y184_I),
.I4(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLM_L_X70Y127_SLICE_X104Y127_CO5),
.O6(CLBLM_L_X70Y127_SLICE_X104Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c393c3c3c6c)
  ) CLBLM_L_X70Y127_SLICE_X104Y127_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(CLBLL_R_X71Y125_SLICE_X106Y125_BO6),
.I2(CLBLM_L_X70Y127_SLICE_X104Y127_AQ),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLM_L_X70Y127_SLICE_X104Y127_CO6),
.O5(CLBLM_L_X70Y127_SLICE_X104Y127_BO5),
.O6(CLBLM_L_X70Y127_SLICE_X104Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00fe11ef0)
  ) CLBLM_L_X70Y127_SLICE_X104Y127_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(CLBLL_R_X73Y122_SLICE_X110Y122_DO6),
.I3(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.I4(CLBLM_L_X70Y128_SLICE_X104Y128_AO6),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_L_X70Y127_SLICE_X104Y127_AO5),
.O6(CLBLM_L_X70Y127_SLICE_X104Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y127_SLICE_X105Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y127_SLICE_X105Y127_DO5),
.O6(CLBLM_L_X70Y127_SLICE_X105Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y127_SLICE_X105Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y127_SLICE_X105Y127_CO5),
.O6(CLBLM_L_X70Y127_SLICE_X105Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y127_SLICE_X105Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y127_SLICE_X105Y127_BO5),
.O6(CLBLM_L_X70Y127_SLICE_X105Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y127_SLICE_X105Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y127_SLICE_X105Y127_AO5),
.O6(CLBLM_L_X70Y127_SLICE_X105Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y128_SLICE_X104Y128_BO6),
.Q(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y128_SLICE_X104Y128_DO5),
.O6(CLBLM_L_X70Y128_SLICE_X104Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y128_SLICE_X104Y128_CO5),
.O6(CLBLM_L_X70Y128_SLICE_X104Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f3f0c0)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_BLUT (
.I0(RIOB33_X105Y181_IOB_X1Y181_I),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I2(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.I3(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I4(CLBLM_L_X70Y127_SLICE_X104Y127_BQ),
.I5(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.O5(CLBLM_L_X70Y128_SLICE_X104Y128_BO5),
.O6(CLBLM_L_X70Y128_SLICE_X104Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1e0f3d1f1e0e2c0)
  ) CLBLM_L_X70Y128_SLICE_X104Y128_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I2(CLBLM_L_X70Y128_SLICE_X104Y128_AQ),
.I3(CLBLM_L_X70Y127_SLICE_X104Y127_BQ),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(RIOB33_X105Y179_IOB_X1Y180_I),
.O5(CLBLM_L_X70Y128_SLICE_X104Y128_AO5),
.O6(CLBLM_L_X70Y128_SLICE_X104Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y128_SLICE_X105Y128_CO6),
.Q(CLBLM_L_X70Y128_SLICE_X105Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y128_SLICE_X105Y128_AO6),
.Q(CLBLM_L_X70Y128_SLICE_X105Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y128_SLICE_X105Y128_DO5),
.O6(CLBLM_L_X70Y128_SLICE_X105Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeff1000fe0010)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_CLUT (
.I0(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I2(CLBLM_L_X70Y128_SLICE_X105Y128_BQ),
.I3(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I4(CLBLM_L_X70Y128_SLICE_X105Y128_AQ),
.I5(RIOB33_X105Y153_IOB_X1Y153_I),
.O5(CLBLM_L_X70Y128_SLICE_X105Y128_CO5),
.O6(CLBLM_L_X70Y128_SLICE_X105Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefdf804040d08)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLM_L_X70Y128_SLICE_X105Y128_BQ),
.I2(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I3(RIOB33_X105Y151_IOB_X1Y152_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(CLBLM_L_X70Y128_SLICE_X105Y128_AQ),
.O5(CLBLM_L_X70Y128_SLICE_X105Y128_BO5),
.O6(CLBLM_L_X70Y128_SLICE_X105Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h666666666666636c)
  ) CLBLM_L_X70Y128_SLICE_X105Y128_ALUT (
.I0(CLBLM_L_X70Y128_SLICE_X105Y128_AQ),
.I1(CLBLL_R_X71Y127_SLICE_X106Y127_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y80_I),
.I3(CLBLM_L_X70Y128_SLICE_X105Y128_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_L_X70Y128_SLICE_X105Y128_AO5),
.O6(CLBLM_L_X70Y128_SLICE_X105Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y129_SLICE_X104Y129_CO6),
.Q(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_L_X70Y129_SLICE_X104Y129_AO6),
.Q(CLBLM_L_X70Y129_SLICE_X104Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y129_SLICE_X104Y129_DO5),
.O6(CLBLM_L_X70Y129_SLICE_X104Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ffe200e2)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_CLUT (
.I0(CLBLM_L_X70Y129_SLICE_X104Y129_BQ),
.I1(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.I2(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I3(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I4(RIOB33_X105Y159_IOB_X1Y159_I),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.O5(CLBLM_L_X70Y129_SLICE_X104Y129_CO5),
.O6(CLBLM_L_X70Y129_SLICE_X104Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0e4f0e4f0ddf088)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLM_L_X70Y129_SLICE_X104Y129_BQ),
.I2(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(RIOB33_X105Y157_IOB_X1Y158_I),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLM_L_X70Y129_SLICE_X104Y129_BO5),
.O6(CLBLM_L_X70Y129_SLICE_X104Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff01de2)
  ) CLBLM_L_X70Y129_SLICE_X104Y129_ALUT (
.I0(CLBLM_L_X70Y129_SLICE_X104Y129_BO6),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLM_L_X70Y129_SLICE_X104Y129_AQ),
.I3(CLBLL_R_X71Y129_SLICE_X106Y129_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y80_I),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLM_L_X70Y129_SLICE_X104Y129_AO5),
.O6(CLBLM_L_X70Y129_SLICE_X104Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y129_SLICE_X105Y129_DO5),
.O6(CLBLM_L_X70Y129_SLICE_X105Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y129_SLICE_X105Y129_CO5),
.O6(CLBLM_L_X70Y129_SLICE_X105Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y129_SLICE_X105Y129_BO5),
.O6(CLBLM_L_X70Y129_SLICE_X105Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X70Y129_SLICE_X105Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X70Y129_SLICE_X105Y129_AO5),
.O6(CLBLM_L_X70Y129_SLICE_X105Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y114_SLICE_X108Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y114_SLICE_X108Y114_DO5),
.O6(CLBLM_L_X72Y114_SLICE_X108Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y114_SLICE_X108Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y114_SLICE_X108Y114_CO5),
.O6(CLBLM_L_X72Y114_SLICE_X108Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y114_SLICE_X108Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y114_SLICE_X108Y114_BO5),
.O6(CLBLM_L_X72Y114_SLICE_X108Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y114_SLICE_X108Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y114_SLICE_X108Y114_AO5),
.O6(CLBLM_L_X72Y114_SLICE_X108Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y114_SLICE_X109Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y114_SLICE_X109Y114_DO5),
.O6(CLBLM_L_X72Y114_SLICE_X109Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fa52d2d5af07878)
  ) CLBLM_L_X72Y114_SLICE_X109Y114_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X72Y115_SLICE_X109Y115_F7BMUX_O),
.I2(CLBLL_R_X71Y119_SLICE_X106Y119_AO6),
.I3(CLBLM_L_X72Y114_SLICE_X109Y114_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_R_X73Y114_SLICE_X110Y114_F8MUX_O),
.O5(CLBLM_L_X72Y114_SLICE_X109Y114_CO5),
.O6(CLBLM_L_X72Y114_SLICE_X109Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cfa0afa0a)
  ) CLBLM_L_X72Y114_SLICE_X109Y114_BLUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I4(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLM_L_X72Y114_SLICE_X109Y114_BO5),
.O6(CLBLM_L_X72Y114_SLICE_X109Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaf0f0cccc)
  ) CLBLM_L_X72Y114_SLICE_X109Y114_ALUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I3(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLM_L_X72Y114_SLICE_X109Y114_AO5),
.O6(CLBLM_L_X72Y114_SLICE_X109Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y114_SLICE_X109Y114_MUXF7A (
.I0(CLBLM_L_X72Y114_SLICE_X109Y114_BO6),
.I1(CLBLM_L_X72Y114_SLICE_X109Y114_AO6),
.O(CLBLM_L_X72Y114_SLICE_X109Y114_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00f0f0aaaa)
  ) CLBLM_L_X72Y115_SLICE_X108Y115_DLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I1(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X72Y115_SLICE_X108Y115_DO5),
.O6(CLBLM_L_X72Y115_SLICE_X108Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88fcfcbb883030)
  ) CLBLM_L_X72Y115_SLICE_X108Y115_CLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.O5(CLBLM_L_X72Y115_SLICE_X108Y115_CO5),
.O6(CLBLM_L_X72Y115_SLICE_X108Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3ee22c0c0ee22)
  ) CLBLM_L_X72Y115_SLICE_X108Y115_BLUT (
.I0(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.O5(CLBLM_L_X72Y115_SLICE_X108Y115_BO5),
.O6(CLBLM_L_X72Y115_SLICE_X108Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccaaaa)
  ) CLBLM_L_X72Y115_SLICE_X108Y115_ALUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I2(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X72Y115_SLICE_X108Y115_AO5),
.O6(CLBLM_L_X72Y115_SLICE_X108Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y115_SLICE_X108Y115_MUXF7A (
.I0(CLBLM_L_X72Y115_SLICE_X108Y115_BO6),
.I1(CLBLM_L_X72Y115_SLICE_X108Y115_AO6),
.O(CLBLM_L_X72Y115_SLICE_X108Y115_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y115_SLICE_X108Y115_MUXF7B (
.I0(CLBLM_L_X72Y115_SLICE_X108Y115_DO6),
.I1(CLBLM_L_X72Y115_SLICE_X108Y115_CO6),
.O(CLBLM_L_X72Y115_SLICE_X108Y115_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X72Y115_SLICE_X108Y115_MUXF8 (
.I0(CLBLM_L_X72Y115_SLICE_X108Y115_F7BMUX_O),
.I1(CLBLM_L_X72Y115_SLICE_X108Y115_F7AMUX_O),
.O(CLBLM_L_X72Y115_SLICE_X108Y115_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cafa0afa0)
  ) CLBLM_L_X72Y115_SLICE_X109Y115_DLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLM_L_X72Y115_SLICE_X109Y115_DO5),
.O6(CLBLM_L_X72Y115_SLICE_X109Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdb97531eca86420)
  ) CLBLM_L_X72Y115_SLICE_X109Y115_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I2(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.O5(CLBLM_L_X72Y115_SLICE_X109Y115_CO5),
.O6(CLBLM_L_X72Y115_SLICE_X109Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fa0afa0a)
  ) CLBLM_L_X72Y115_SLICE_X109Y115_BLUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I4(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X72Y115_SLICE_X109Y115_BO5),
.O6(CLBLM_L_X72Y115_SLICE_X109Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0acfcffa0ac0c0)
  ) CLBLM_L_X72Y115_SLICE_X109Y115_ALUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.O5(CLBLM_L_X72Y115_SLICE_X109Y115_AO5),
.O6(CLBLM_L_X72Y115_SLICE_X109Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y115_SLICE_X109Y115_MUXF7A (
.I0(CLBLM_L_X72Y115_SLICE_X109Y115_BO6),
.I1(CLBLM_L_X72Y115_SLICE_X109Y115_AO6),
.O(CLBLM_L_X72Y115_SLICE_X109Y115_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y115_SLICE_X109Y115_MUXF7B (
.I0(CLBLM_L_X72Y115_SLICE_X109Y115_DO6),
.I1(CLBLM_L_X72Y115_SLICE_X109Y115_CO6),
.O(CLBLM_L_X72Y115_SLICE_X109Y115_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h666633cc3c3c3c3c)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_DLUT (
.I0(CLBLM_L_X72Y117_SLICE_X108Y117_F7BMUX_O),
.I1(CLBLM_L_X70Y124_SLICE_X104Y124_CO6),
.I2(CLBLM_L_X72Y115_SLICE_X108Y115_F8MUX_O),
.I3(CLBLM_L_X72Y116_SLICE_X108Y116_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLM_L_X72Y116_SLICE_X108Y116_DO5),
.O6(CLBLM_L_X72Y116_SLICE_X108Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h56a656a65555aaaa)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_CLUT (
.I0(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.I1(CLBLM_L_X72Y116_SLICE_X109Y116_F7AMUX_O),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(CLBLM_L_X72Y117_SLICE_X108Y117_F7AMUX_O),
.I4(CLBLM_L_X74Y116_SLICE_X112Y116_F8MUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLM_L_X72Y116_SLICE_X108Y116_CO5),
.O6(CLBLM_L_X72Y116_SLICE_X108Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cfcfafa0c0c0)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_BLUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.O5(CLBLM_L_X72Y116_SLICE_X108Y116_BO5),
.O6(CLBLM_L_X72Y116_SLICE_X108Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0acfcffa0ac0c0)
  ) CLBLM_L_X72Y116_SLICE_X108Y116_ALUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.O5(CLBLM_L_X72Y116_SLICE_X108Y116_AO5),
.O6(CLBLM_L_X72Y116_SLICE_X108Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y116_SLICE_X108Y116_MUXF7A (
.I0(CLBLM_L_X72Y116_SLICE_X108Y116_BO6),
.I1(CLBLM_L_X72Y116_SLICE_X108Y116_AO6),
.O(CLBLM_L_X72Y116_SLICE_X108Y116_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heef322f3eec022c0)
  ) CLBLM_L_X72Y116_SLICE_X109Y116_DLUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLM_L_X72Y116_SLICE_X109Y116_DO5),
.O6(CLBLM_L_X72Y116_SLICE_X109Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcaffca00caf0ca0)
  ) CLBLM_L_X72Y116_SLICE_X109Y116_CLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I1(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.O5(CLBLM_L_X72Y116_SLICE_X109Y116_CO5),
.O6(CLBLM_L_X72Y116_SLICE_X109Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe5eae04f454a40)
  ) CLBLM_L_X72Y116_SLICE_X109Y116_BLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.O5(CLBLM_L_X72Y116_SLICE_X109Y116_BO5),
.O6(CLBLM_L_X72Y116_SLICE_X109Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0fcfcafa00c0c)
  ) CLBLM_L_X72Y116_SLICE_X109Y116_ALUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.O5(CLBLM_L_X72Y116_SLICE_X109Y116_AO5),
.O6(CLBLM_L_X72Y116_SLICE_X109Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y116_SLICE_X109Y116_MUXF7A (
.I0(CLBLM_L_X72Y116_SLICE_X109Y116_BO6),
.I1(CLBLM_L_X72Y116_SLICE_X109Y116_AO6),
.O(CLBLM_L_X72Y116_SLICE_X109Y116_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y116_SLICE_X109Y116_MUXF7B (
.I0(CLBLM_L_X72Y116_SLICE_X109Y116_DO6),
.I1(CLBLM_L_X72Y116_SLICE_X109Y116_CO6),
.O(CLBLM_L_X72Y116_SLICE_X109Y116_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fafa0a0a)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_DLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X72Y117_SLICE_X108Y117_DO5),
.O6(CLBLM_L_X72Y117_SLICE_X108Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef2cec23e320e02)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_CLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.O5(CLBLM_L_X72Y117_SLICE_X108Y117_CO5),
.O6(CLBLM_L_X72Y117_SLICE_X108Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0caca0f00caca)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_BLUT (
.I0(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.O5(CLBLM_L_X72Y117_SLICE_X108Y117_BO5),
.O6(CLBLM_L_X72Y117_SLICE_X108Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbcbf8c83b0b3808)
  ) CLBLM_L_X72Y117_SLICE_X108Y117_ALUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I4(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLM_L_X72Y117_SLICE_X108Y117_AO5),
.O6(CLBLM_L_X72Y117_SLICE_X108Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y117_SLICE_X108Y117_MUXF7A (
.I0(CLBLM_L_X72Y117_SLICE_X108Y117_BO6),
.I1(CLBLM_L_X72Y117_SLICE_X108Y117_AO6),
.O(CLBLM_L_X72Y117_SLICE_X108Y117_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y117_SLICE_X108Y117_MUXF7B (
.I0(CLBLM_L_X72Y117_SLICE_X108Y117_DO6),
.I1(CLBLM_L_X72Y117_SLICE_X108Y117_CO6),
.O(CLBLM_L_X72Y117_SLICE_X108Y117_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X109Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X109Y117_DO5),
.O6(CLBLM_L_X72Y117_SLICE_X109Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y117_SLICE_X109Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y117_SLICE_X109Y117_CO5),
.O6(CLBLM_L_X72Y117_SLICE_X109Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfa0cfafc0a0c0a)
  ) CLBLM_L_X72Y117_SLICE_X109Y117_BLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.O5(CLBLM_L_X72Y117_SLICE_X109Y117_BO5),
.O6(CLBLM_L_X72Y117_SLICE_X109Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcaf0caffca00ca0)
  ) CLBLM_L_X72Y117_SLICE_X109Y117_ALUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLM_L_X72Y117_SLICE_X109Y117_AO5),
.O6(CLBLM_L_X72Y117_SLICE_X109Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y117_SLICE_X109Y117_MUXF7A (
.I0(CLBLM_L_X72Y117_SLICE_X109Y117_BO6),
.I1(CLBLM_L_X72Y117_SLICE_X109Y117_AO6),
.O(CLBLM_L_X72Y117_SLICE_X109Y117_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1b1be4e411bbee44)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_DLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLL_R_X73Y118_SLICE_X110Y118_F8MUX_O),
.I2(CLBLM_L_X72Y118_SLICE_X109Y118_F7BMUX_O),
.I3(CLBLM_L_X72Y118_SLICE_X108Y118_F7AMUX_O),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_DO6),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_L_X72Y118_SLICE_X108Y118_DO5),
.O6(CLBLM_L_X72Y118_SLICE_X108Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h02a2fd5d57f7a808)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X72Y118_SLICE_X109Y118_F7AMUX_O),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(CLBLM_L_X72Y117_SLICE_X109Y117_F7AMUX_O),
.I4(CLBLM_L_X70Y119_SLICE_X105Y119_CO6),
.I5(CLBLL_R_X71Y118_SLICE_X107Y118_F8MUX_O),
.O5(CLBLM_L_X72Y118_SLICE_X108Y118_CO5),
.O6(CLBLM_L_X72Y118_SLICE_X108Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaaffaa00)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_BLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I1(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLM_L_X72Y118_SLICE_X108Y118_BO5),
.O6(CLBLM_L_X72Y118_SLICE_X108Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cfcfc0c0)
  ) CLBLM_L_X72Y118_SLICE_X108Y118_ALUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLM_L_X72Y118_SLICE_X108Y118_AO5),
.O6(CLBLM_L_X72Y118_SLICE_X108Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y118_SLICE_X108Y118_MUXF7A (
.I0(CLBLM_L_X72Y118_SLICE_X108Y118_BO6),
.I1(CLBLM_L_X72Y118_SLICE_X108Y118_AO6),
.O(CLBLM_L_X72Y118_SLICE_X108Y118_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdecb9a875643120)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_DLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.O5(CLBLM_L_X72Y118_SLICE_X109Y118_DO5),
.O6(CLBLM_L_X72Y118_SLICE_X109Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heefaee5044fa4450)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.O5(CLBLM_L_X72Y118_SLICE_X109Y118_CO5),
.O6(CLBLM_L_X72Y118_SLICE_X109Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55d8d8aa00d8d8)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.O5(CLBLM_L_X72Y118_SLICE_X109Y118_BO5),
.O6(CLBLM_L_X72Y118_SLICE_X109Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fcacaf000caca)
  ) CLBLM_L_X72Y118_SLICE_X109Y118_ALUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I1(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.O5(CLBLM_L_X72Y118_SLICE_X109Y118_AO5),
.O6(CLBLM_L_X72Y118_SLICE_X109Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y118_SLICE_X109Y118_MUXF7A (
.I0(CLBLM_L_X72Y118_SLICE_X109Y118_BO6),
.I1(CLBLM_L_X72Y118_SLICE_X109Y118_AO6),
.O(CLBLM_L_X72Y118_SLICE_X109Y118_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y118_SLICE_X109Y118_MUXF7B (
.I0(CLBLM_L_X72Y118_SLICE_X109Y118_DO6),
.I1(CLBLM_L_X72Y118_SLICE_X109Y118_CO6),
.O(CLBLM_L_X72Y118_SLICE_X109Y118_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h220a775fddf588a0)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_DLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X72Y119_SLICE_X109Y119_F7BMUX_O),
.I2(CLBLL_R_X71Y119_SLICE_X107Y119_F7AMUX_O),
.I3(LIOB33_X0Y81_IOB_X0Y81_I),
.I4(CLBLM_L_X72Y121_SLICE_X108Y121_F8MUX_O),
.I5(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.O5(CLBLM_L_X72Y119_SLICE_X108Y119_DO5),
.O6(CLBLM_L_X72Y119_SLICE_X108Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2727d8d805affa50)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X72Y119_SLICE_X109Y119_F7AMUX_O),
.I2(CLBLL_R_X73Y119_SLICE_X110Y119_F8MUX_O),
.I3(CLBLM_L_X72Y119_SLICE_X108Y119_F7AMUX_O),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_DO6),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_L_X72Y119_SLICE_X108Y119_CO5),
.O6(CLBLM_L_X72Y119_SLICE_X108Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb3bcb0bf838c808)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_BLUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I4(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.O5(CLBLM_L_X72Y119_SLICE_X108Y119_BO5),
.O6(CLBLM_L_X72Y119_SLICE_X108Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfafcfa0c0afc0a0)
  ) CLBLM_L_X72Y119_SLICE_X108Y119_ALUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I5(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.O5(CLBLM_L_X72Y119_SLICE_X108Y119_AO5),
.O6(CLBLM_L_X72Y119_SLICE_X108Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y119_SLICE_X108Y119_MUXF7A (
.I0(CLBLM_L_X72Y119_SLICE_X108Y119_BO6),
.I1(CLBLM_L_X72Y119_SLICE_X108Y119_AO6),
.O(CLBLM_L_X72Y119_SLICE_X108Y119_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_DLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X72Y119_SLICE_X109Y119_DO5),
.O6(CLBLM_L_X72Y119_SLICE_X109Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_CLUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I2(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X72Y119_SLICE_X109Y119_CO5),
.O6(CLBLM_L_X72Y119_SLICE_X109Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcbb883030bb88)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_BLUT (
.I0(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.O5(CLBLM_L_X72Y119_SLICE_X109Y119_BO5),
.O6(CLBLM_L_X72Y119_SLICE_X109Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffac0facf0ac00ac)
  ) CLBLM_L_X72Y119_SLICE_X109Y119_ALUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.O5(CLBLM_L_X72Y119_SLICE_X109Y119_AO5),
.O6(CLBLM_L_X72Y119_SLICE_X109Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y119_SLICE_X109Y119_MUXF7A (
.I0(CLBLM_L_X72Y119_SLICE_X109Y119_BO6),
.I1(CLBLM_L_X72Y119_SLICE_X109Y119_AO6),
.O(CLBLM_L_X72Y119_SLICE_X109Y119_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y119_SLICE_X109Y119_MUXF7B (
.I0(CLBLM_L_X72Y119_SLICE_X109Y119_DO6),
.I1(CLBLM_L_X72Y119_SLICE_X109Y119_CO6),
.O(CLBLM_L_X72Y119_SLICE_X109Y119_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h339366c639996ccc)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_DLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X70Y119_SLICE_X105Y119_CO6),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(CLBLM_L_X72Y120_SLICE_X108Y120_F7AMUX_O),
.I4(CLBLM_L_X72Y121_SLICE_X109Y121_F8MUX_O),
.I5(CLBLL_R_X71Y120_SLICE_X106Y120_F7BMUX_O),
.O5(CLBLM_L_X72Y120_SLICE_X108Y120_DO5),
.O6(CLBLM_L_X72Y120_SLICE_X108Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd32c8c6778961de1)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_CLUT (
.I0(CLBLL_R_X71Y122_SLICE_X106Y122_AO6),
.I1(CLBLM_L_X74Y120_SLICE_X113Y120_AO6),
.I2(CLBLL_R_X71Y120_SLICE_X107Y120_AO6),
.I3(CLBLL_R_X73Y120_SLICE_X111Y120_DO6),
.I4(CLBLM_L_X72Y120_SLICE_X108Y120_DO6),
.I5(CLBLL_R_X73Y120_SLICE_X111Y120_CO6),
.O5(CLBLM_L_X72Y120_SLICE_X108Y120_CO5),
.O6(CLBLM_L_X72Y120_SLICE_X108Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_BLUT (
.I0(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I3(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y120_SLICE_X108Y120_BO5),
.O6(CLBLM_L_X72Y120_SLICE_X108Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccff00aaaa)
  ) CLBLM_L_X72Y120_SLICE_X108Y120_ALUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y120_SLICE_X108Y120_AO5),
.O6(CLBLM_L_X72Y120_SLICE_X108Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y120_SLICE_X108Y120_MUXF7A (
.I0(CLBLM_L_X72Y120_SLICE_X108Y120_BO6),
.I1(CLBLM_L_X72Y120_SLICE_X108Y120_AO6),
.O(CLBLM_L_X72Y120_SLICE_X108Y120_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ffd855d8aad800)
  ) CLBLM_L_X72Y120_SLICE_X109Y120_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.O5(CLBLM_L_X72Y120_SLICE_X109Y120_DO5),
.O6(CLBLM_L_X72Y120_SLICE_X109Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0aacc00f0aacc)
  ) CLBLM_L_X72Y120_SLICE_X109Y120_CLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.O5(CLBLM_L_X72Y120_SLICE_X109Y120_CO5),
.O6(CLBLM_L_X72Y120_SLICE_X109Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLM_L_X72Y120_SLICE_X109Y120_BLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I1(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y120_SLICE_X109Y120_BO5),
.O6(CLBLM_L_X72Y120_SLICE_X109Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55d8d8aa00d8d8)
  ) CLBLM_L_X72Y120_SLICE_X109Y120_ALUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.O5(CLBLM_L_X72Y120_SLICE_X109Y120_AO5),
.O6(CLBLM_L_X72Y120_SLICE_X109Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y120_SLICE_X109Y120_MUXF7A (
.I0(CLBLM_L_X72Y120_SLICE_X109Y120_BO6),
.I1(CLBLM_L_X72Y120_SLICE_X109Y120_AO6),
.O(CLBLM_L_X72Y120_SLICE_X109Y120_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y120_SLICE_X109Y120_MUXF7B (
.I0(CLBLM_L_X72Y120_SLICE_X109Y120_DO6),
.I1(CLBLM_L_X72Y120_SLICE_X109Y120_CO6),
.O(CLBLM_L_X72Y120_SLICE_X109Y120_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X72Y120_SLICE_X109Y120_MUXF8 (
.I0(CLBLM_L_X72Y120_SLICE_X109Y120_F7BMUX_O),
.I1(CLBLM_L_X72Y120_SLICE_X109Y120_F7AMUX_O),
.O(CLBLM_L_X72Y120_SLICE_X109Y120_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee50eefa445044)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_DLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.O5(CLBLM_L_X72Y121_SLICE_X108Y121_DO5),
.O6(CLBLM_L_X72Y121_SLICE_X108Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5eea0eef544a044)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_CLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I5(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.O5(CLBLM_L_X72Y121_SLICE_X108Y121_CO5),
.O6(CLBLM_L_X72Y121_SLICE_X108Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2ffcce2e23300)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_BLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I3(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.O5(CLBLM_L_X72Y121_SLICE_X108Y121_BO5),
.O6(CLBLM_L_X72Y121_SLICE_X108Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300e2e2e2e2)
  ) CLBLM_L_X72Y121_SLICE_X108Y121_ALUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y121_SLICE_X108Y121_AO5),
.O6(CLBLM_L_X72Y121_SLICE_X108Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y121_SLICE_X108Y121_MUXF7A (
.I0(CLBLM_L_X72Y121_SLICE_X108Y121_BO6),
.I1(CLBLM_L_X72Y121_SLICE_X108Y121_AO6),
.O(CLBLM_L_X72Y121_SLICE_X108Y121_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y121_SLICE_X108Y121_MUXF7B (
.I0(CLBLM_L_X72Y121_SLICE_X108Y121_DO6),
.I1(CLBLM_L_X72Y121_SLICE_X108Y121_CO6),
.O(CLBLM_L_X72Y121_SLICE_X108Y121_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X72Y121_SLICE_X108Y121_MUXF8 (
.I0(CLBLM_L_X72Y121_SLICE_X108Y121_F7BMUX_O),
.I1(CLBLM_L_X72Y121_SLICE_X108Y121_F7AMUX_O),
.O(CLBLM_L_X72Y121_SLICE_X108Y121_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe3ece02f232c20)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_DLUT (
.I0(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.O5(CLBLM_L_X72Y121_SLICE_X109Y121_DO5),
.O6(CLBLM_L_X72Y121_SLICE_X109Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2ffcce2e23300)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_CLUT (
.I0(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I3(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.O5(CLBLM_L_X72Y121_SLICE_X109Y121_CO5),
.O6(CLBLM_L_X72Y121_SLICE_X109Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50eeee4444)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_BLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I2(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y121_SLICE_X109Y121_BO5),
.O6(CLBLM_L_X72Y121_SLICE_X109Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5dd88a0a0dd88)
  ) CLBLM_L_X72Y121_SLICE_X109Y121_ALUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.O5(CLBLM_L_X72Y121_SLICE_X109Y121_AO5),
.O6(CLBLM_L_X72Y121_SLICE_X109Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y121_SLICE_X109Y121_MUXF7A (
.I0(CLBLM_L_X72Y121_SLICE_X109Y121_BO6),
.I1(CLBLM_L_X72Y121_SLICE_X109Y121_AO6),
.O(CLBLM_L_X72Y121_SLICE_X109Y121_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y121_SLICE_X109Y121_MUXF7B (
.I0(CLBLM_L_X72Y121_SLICE_X109Y121_DO6),
.I1(CLBLM_L_X72Y121_SLICE_X109Y121_CO6),
.O(CLBLM_L_X72Y121_SLICE_X109Y121_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X72Y121_SLICE_X109Y121_MUXF8 (
.I0(CLBLM_L_X72Y121_SLICE_X109Y121_F7BMUX_O),
.I1(CLBLM_L_X72Y121_SLICE_X109Y121_F7AMUX_O),
.O(CLBLM_L_X72Y121_SLICE_X109Y121_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X108Y122_DO5),
.O6(CLBLM_L_X72Y122_SLICE_X108Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X108Y122_CO5),
.O6(CLBLM_L_X72Y122_SLICE_X108Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X108Y122_BO5),
.O6(CLBLM_L_X72Y122_SLICE_X108Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33c366663ccc6666)
  ) CLBLM_L_X72Y122_SLICE_X108Y122_ALUT (
.I0(CLBLM_L_X72Y123_SLICE_X109Y123_F8MUX_O),
.I1(CLBLL_L_X2Y120_SLICE_X0Y120_DO6),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(CLBLM_L_X72Y123_SLICE_X108Y123_F7BMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLM_L_X72Y123_SLICE_X108Y123_F7AMUX_O),
.O5(CLBLM_L_X72Y122_SLICE_X108Y122_AO5),
.O6(CLBLM_L_X72Y122_SLICE_X108Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X109Y122_DO5),
.O6(CLBLM_L_X72Y122_SLICE_X109Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X109Y122_CO5),
.O6(CLBLM_L_X72Y122_SLICE_X109Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X109Y122_BO5),
.O6(CLBLM_L_X72Y122_SLICE_X109Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y122_SLICE_X109Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y122_SLICE_X109Y122_AO5),
.O6(CLBLM_L_X72Y122_SLICE_X109Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfc0cfc0)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_DLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I4(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y123_SLICE_X108Y123_DO5),
.O6(CLBLM_L_X72Y123_SLICE_X108Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfa0cfafc0a0c0a)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_CLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I5(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.O5(CLBLM_L_X72Y123_SLICE_X108Y123_CO5),
.O6(CLBLM_L_X72Y123_SLICE_X108Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0ee44ee44)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_BLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I2(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y123_SLICE_X108Y123_BO5),
.O6(CLBLM_L_X72Y123_SLICE_X108Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ffcc3300)
  ) CLBLM_L_X72Y123_SLICE_X108Y123_ALUT (
.I0(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I4(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y123_SLICE_X108Y123_AO5),
.O6(CLBLM_L_X72Y123_SLICE_X108Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y123_SLICE_X108Y123_MUXF7A (
.I0(CLBLM_L_X72Y123_SLICE_X108Y123_BO6),
.I1(CLBLM_L_X72Y123_SLICE_X108Y123_AO6),
.O(CLBLM_L_X72Y123_SLICE_X108Y123_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y123_SLICE_X108Y123_MUXF7B (
.I0(CLBLM_L_X72Y123_SLICE_X108Y123_DO6),
.I1(CLBLM_L_X72Y123_SLICE_X108Y123_CO6),
.O(CLBLM_L_X72Y123_SLICE_X108Y123_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf8fbc8cb383b080)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_DLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I5(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.O5(CLBLM_L_X72Y123_SLICE_X109Y123_DO5),
.O6(CLBLM_L_X72Y123_SLICE_X109Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef23e32cec20e02)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_CLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I5(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.O5(CLBLM_L_X72Y123_SLICE_X109Y123_CO5),
.O6(CLBLM_L_X72Y123_SLICE_X109Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ff55aa00)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_BLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I2(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y123_SLICE_X109Y123_BO5),
.O6(CLBLM_L_X72Y123_SLICE_X109Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44f5f5a0a0)
  ) CLBLM_L_X72Y123_SLICE_X109Y123_ALUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I4(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y123_SLICE_X109Y123_AO5),
.O6(CLBLM_L_X72Y123_SLICE_X109Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y123_SLICE_X109Y123_MUXF7A (
.I0(CLBLM_L_X72Y123_SLICE_X109Y123_BO6),
.I1(CLBLM_L_X72Y123_SLICE_X109Y123_AO6),
.O(CLBLM_L_X72Y123_SLICE_X109Y123_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y123_SLICE_X109Y123_MUXF7B (
.I0(CLBLM_L_X72Y123_SLICE_X109Y123_DO6),
.I1(CLBLM_L_X72Y123_SLICE_X109Y123_CO6),
.O(CLBLM_L_X72Y123_SLICE_X109Y123_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X72Y123_SLICE_X109Y123_MUXF8 (
.I0(CLBLM_L_X72Y123_SLICE_X109Y123_F7BMUX_O),
.I1(CLBLM_L_X72Y123_SLICE_X109Y123_F7AMUX_O),
.O(CLBLM_L_X72Y123_SLICE_X109Y123_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y124_SLICE_X108Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y124_SLICE_X108Y124_DO5),
.O6(CLBLM_L_X72Y124_SLICE_X108Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a555aaa665566aa)
  ) CLBLM_L_X72Y124_SLICE_X108Y124_CLUT (
.I0(CLBLM_L_X70Y123_SLICE_X104Y123_BO6),
.I1(CLBLM_L_X72Y124_SLICE_X109Y124_F7AMUX_O),
.I2(CLBLM_L_X72Y124_SLICE_X109Y124_F7BMUX_O),
.I3(LIOB33_X0Y81_IOB_X0Y82_I),
.I4(CLBLL_R_X73Y124_SLICE_X110Y124_F8MUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_L_X72Y124_SLICE_X108Y124_CO5),
.O6(CLBLM_L_X72Y124_SLICE_X108Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef2fe323ec2ce020)
  ) CLBLM_L_X72Y124_SLICE_X108Y124_BLUT (
.I0(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I5(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.O5(CLBLM_L_X72Y124_SLICE_X108Y124_BO5),
.O6(CLBLM_L_X72Y124_SLICE_X108Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf8fda8ad585d080)
  ) CLBLM_L_X72Y124_SLICE_X108Y124_ALUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.O5(CLBLM_L_X72Y124_SLICE_X108Y124_AO5),
.O6(CLBLM_L_X72Y124_SLICE_X108Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y124_SLICE_X108Y124_MUXF7A (
.I0(CLBLM_L_X72Y124_SLICE_X108Y124_BO6),
.I1(CLBLM_L_X72Y124_SLICE_X108Y124_AO6),
.O(CLBLM_L_X72Y124_SLICE_X108Y124_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLM_L_X72Y124_SLICE_X109Y124_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I2(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I4(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y124_SLICE_X109Y124_DO5),
.O6(CLBLM_L_X72Y124_SLICE_X109Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccaaaaff00)
  ) CLBLM_L_X72Y124_SLICE_X109Y124_CLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y124_SLICE_X109Y124_CO5),
.O6(CLBLM_L_X72Y124_SLICE_X109Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0ddddf5a08888)
  ) CLBLM_L_X72Y124_SLICE_X109Y124_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I2(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.O5(CLBLM_L_X72Y124_SLICE_X109Y124_BO5),
.O6(CLBLM_L_X72Y124_SLICE_X109Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaafff0ccaa00f0)
  ) CLBLM_L_X72Y124_SLICE_X109Y124_ALUT (
.I0(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.O5(CLBLM_L_X72Y124_SLICE_X109Y124_AO5),
.O6(CLBLM_L_X72Y124_SLICE_X109Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y124_SLICE_X109Y124_MUXF7A (
.I0(CLBLM_L_X72Y124_SLICE_X109Y124_BO6),
.I1(CLBLM_L_X72Y124_SLICE_X109Y124_AO6),
.O(CLBLM_L_X72Y124_SLICE_X109Y124_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y124_SLICE_X109Y124_MUXF7B (
.I0(CLBLM_L_X72Y124_SLICE_X109Y124_DO6),
.I1(CLBLM_L_X72Y124_SLICE_X109Y124_CO6),
.O(CLBLM_L_X72Y124_SLICE_X109Y124_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbd9eac873516240)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.O5(CLBLM_L_X72Y125_SLICE_X108Y125_DO5),
.O6(CLBLM_L_X72Y125_SLICE_X108Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdadf8a85d0d5808)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I5(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.O5(CLBLM_L_X72Y125_SLICE_X108Y125_CO5),
.O6(CLBLM_L_X72Y125_SLICE_X108Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0aaccaacc)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_BLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y125_SLICE_X108Y125_BO5),
.O6(CLBLM_L_X72Y125_SLICE_X108Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaef4a45e0e5404)
  ) CLBLM_L_X72Y125_SLICE_X108Y125_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.O5(CLBLM_L_X72Y125_SLICE_X108Y125_AO5),
.O6(CLBLM_L_X72Y125_SLICE_X108Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y125_SLICE_X108Y125_MUXF7A (
.I0(CLBLM_L_X72Y125_SLICE_X108Y125_BO6),
.I1(CLBLM_L_X72Y125_SLICE_X108Y125_AO6),
.O(CLBLM_L_X72Y125_SLICE_X108Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y125_SLICE_X108Y125_MUXF7B (
.I0(CLBLM_L_X72Y125_SLICE_X108Y125_DO6),
.I1(CLBLM_L_X72Y125_SLICE_X108Y125_CO6),
.O(CLBLM_L_X72Y125_SLICE_X108Y125_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_DLUT (
.I0(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I2(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y125_SLICE_X109Y125_DO5),
.O6(CLBLM_L_X72Y125_SLICE_X109Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafcfa0c0afc0a0c)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_CLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.O5(CLBLM_L_X72Y125_SLICE_X109Y125_CO5),
.O6(CLBLM_L_X72Y125_SLICE_X109Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdad5d08f8a8580)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_BLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.O5(CLBLM_L_X72Y125_SLICE_X109Y125_BO5),
.O6(CLBLM_L_X72Y125_SLICE_X109Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5eea0eef544a044)
  ) CLBLM_L_X72Y125_SLICE_X109Y125_ALUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.O5(CLBLM_L_X72Y125_SLICE_X109Y125_AO5),
.O6(CLBLM_L_X72Y125_SLICE_X109Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y125_SLICE_X109Y125_MUXF7A (
.I0(CLBLM_L_X72Y125_SLICE_X109Y125_BO6),
.I1(CLBLM_L_X72Y125_SLICE_X109Y125_AO6),
.O(CLBLM_L_X72Y125_SLICE_X109Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y125_SLICE_X109Y125_MUXF7B (
.I0(CLBLM_L_X72Y125_SLICE_X109Y125_DO6),
.I1(CLBLM_L_X72Y125_SLICE_X109Y125_CO6),
.O(CLBLM_L_X72Y125_SLICE_X109Y125_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X72Y125_SLICE_X109Y125_MUXF8 (
.I0(CLBLM_L_X72Y125_SLICE_X109Y125_F7BMUX_O),
.I1(CLBLM_L_X72Y125_SLICE_X109Y125_F7AMUX_O),
.O(CLBLM_L_X72Y125_SLICE_X109Y125_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5eef544a0eea044)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I2(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.O5(CLBLM_L_X72Y126_SLICE_X108Y126_DO5),
.O6(CLBLM_L_X72Y126_SLICE_X108Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccffaaf0cc00aa)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_CLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I2(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.O5(CLBLM_L_X72Y126_SLICE_X108Y126_CO5),
.O6(CLBLM_L_X72Y126_SLICE_X108Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30bbbb8888)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_BLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y126_SLICE_X108Y126_BO5),
.O6(CLBLM_L_X72Y126_SLICE_X108Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00f0f0aaaa)
  ) CLBLM_L_X72Y126_SLICE_X108Y126_ALUT (
.I0(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I2(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y126_SLICE_X108Y126_AO5),
.O6(CLBLM_L_X72Y126_SLICE_X108Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y126_SLICE_X108Y126_MUXF7A (
.I0(CLBLM_L_X72Y126_SLICE_X108Y126_BO6),
.I1(CLBLM_L_X72Y126_SLICE_X108Y126_AO6),
.O(CLBLM_L_X72Y126_SLICE_X108Y126_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y126_SLICE_X108Y126_MUXF7B (
.I0(CLBLM_L_X72Y126_SLICE_X108Y126_DO6),
.I1(CLBLM_L_X72Y126_SLICE_X108Y126_CO6),
.O(CLBLM_L_X72Y126_SLICE_X108Y126_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X72Y126_SLICE_X108Y126_MUXF8 (
.I0(CLBLM_L_X72Y126_SLICE_X108Y126_F7BMUX_O),
.I1(CLBLM_L_X72Y126_SLICE_X108Y126_F7AMUX_O),
.O(CLBLM_L_X72Y126_SLICE_X108Y126_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbcb3b0bf8c83808)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_DLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I4(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I5(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.O5(CLBLM_L_X72Y126_SLICE_X109Y126_DO5),
.O6(CLBLM_L_X72Y126_SLICE_X109Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee50eefa445044)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I2(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.O5(CLBLM_L_X72Y126_SLICE_X109Y126_CO5),
.O6(CLBLM_L_X72Y126_SLICE_X109Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888f3c0f3c0)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_BLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y126_SLICE_X109Y126_BO5),
.O6(CLBLM_L_X72Y126_SLICE_X109Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLM_L_X72Y126_SLICE_X109Y126_ALUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y126_SLICE_X109Y126_AO5),
.O6(CLBLM_L_X72Y126_SLICE_X109Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y126_SLICE_X109Y126_MUXF7A (
.I0(CLBLM_L_X72Y126_SLICE_X109Y126_BO6),
.I1(CLBLM_L_X72Y126_SLICE_X109Y126_AO6),
.O(CLBLM_L_X72Y126_SLICE_X109Y126_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y126_SLICE_X109Y126_MUXF7B (
.I0(CLBLM_L_X72Y126_SLICE_X109Y126_DO6),
.I1(CLBLM_L_X72Y126_SLICE_X109Y126_CO6),
.O(CLBLM_L_X72Y126_SLICE_X109Y126_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefea4f4ae5e04540)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.O5(CLBLM_L_X72Y127_SLICE_X108Y127_DO5),
.O6(CLBLM_L_X72Y127_SLICE_X108Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf8fda8ad585d080)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.O5(CLBLM_L_X72Y127_SLICE_X108Y127_CO5),
.O6(CLBLM_L_X72Y127_SLICE_X108Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_BLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y127_SLICE_X108Y127_BO5),
.O6(CLBLM_L_X72Y127_SLICE_X108Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0acfcffa0ac0c0)
  ) CLBLM_L_X72Y127_SLICE_X108Y127_ALUT (
.I0(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I1(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.O5(CLBLM_L_X72Y127_SLICE_X108Y127_AO5),
.O6(CLBLM_L_X72Y127_SLICE_X108Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y127_SLICE_X108Y127_MUXF7A (
.I0(CLBLM_L_X72Y127_SLICE_X108Y127_BO6),
.I1(CLBLM_L_X72Y127_SLICE_X108Y127_AO6),
.O(CLBLM_L_X72Y127_SLICE_X108Y127_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y127_SLICE_X108Y127_MUXF7B (
.I0(CLBLM_L_X72Y127_SLICE_X108Y127_DO6),
.I1(CLBLM_L_X72Y127_SLICE_X108Y127_CO6),
.O(CLBLM_L_X72Y127_SLICE_X108Y127_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ffaa5500)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y127_SLICE_X109Y127_DO5),
.O6(CLBLM_L_X72Y127_SLICE_X109Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fafa5050)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I2(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y127_SLICE_X109Y127_CO5),
.O6(CLBLM_L_X72Y127_SLICE_X109Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe5eae0ef454a404)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_BLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I5(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.O5(CLBLM_L_X72Y127_SLICE_X109Y127_BO5),
.O6(CLBLM_L_X72Y127_SLICE_X109Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cfcfafa0c0c0)
  ) CLBLM_L_X72Y127_SLICE_X109Y127_ALUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.O5(CLBLM_L_X72Y127_SLICE_X109Y127_AO5),
.O6(CLBLM_L_X72Y127_SLICE_X109Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y127_SLICE_X109Y127_MUXF7A (
.I0(CLBLM_L_X72Y127_SLICE_X109Y127_BO6),
.I1(CLBLM_L_X72Y127_SLICE_X109Y127_AO6),
.O(CLBLM_L_X72Y127_SLICE_X109Y127_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y127_SLICE_X109Y127_MUXF7B (
.I0(CLBLM_L_X72Y127_SLICE_X109Y127_DO6),
.I1(CLBLM_L_X72Y127_SLICE_X109Y127_CO6),
.O(CLBLM_L_X72Y127_SLICE_X109Y127_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X72Y127_SLICE_X109Y127_MUXF8 (
.I0(CLBLM_L_X72Y127_SLICE_X109Y127_F7BMUX_O),
.I1(CLBLM_L_X72Y127_SLICE_X109Y127_F7AMUX_O),
.O(CLBLM_L_X72Y127_SLICE_X109Y127_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y128_SLICE_X108Y128_DO5),
.O6(CLBLM_L_X72Y128_SLICE_X108Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h369c369c36369c9c)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLL_R_X71Y131_SLICE_X106Y131_CO6),
.I2(CLBLM_L_X72Y129_SLICE_X108Y129_F8MUX_O),
.I3(CLBLM_L_X72Y128_SLICE_X108Y128_F7AMUX_O),
.I4(CLBLM_L_X72Y129_SLICE_X109Y129_F7AMUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_L_X72Y128_SLICE_X108Y128_CO5),
.O6(CLBLM_L_X72Y128_SLICE_X108Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfa0cfafc0a0c0a)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_BLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.O5(CLBLM_L_X72Y128_SLICE_X108Y128_BO5),
.O6(CLBLM_L_X72Y128_SLICE_X108Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe5ef454ae0ea404)
  ) CLBLM_L_X72Y128_SLICE_X108Y128_ALUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.O5(CLBLM_L_X72Y128_SLICE_X108Y128_AO5),
.O6(CLBLM_L_X72Y128_SLICE_X108Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y128_SLICE_X108Y128_MUXF7A (
.I0(CLBLM_L_X72Y128_SLICE_X108Y128_BO6),
.I1(CLBLM_L_X72Y128_SLICE_X108Y128_AO6),
.O(CLBLM_L_X72Y128_SLICE_X108Y128_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h440fbbf0770f88f0)
  ) CLBLM_L_X72Y128_SLICE_X109Y128_DLUT (
.I0(CLBLM_L_X72Y129_SLICE_X109Y129_F7BMUX_O),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLM_L_X74Y128_SLICE_X113Y128_F8MUX_O),
.I3(LIOB33_X0Y81_IOB_X0Y82_I),
.I4(CLBLM_L_X70Y128_SLICE_X104Y128_BO6),
.I5(CLBLL_R_X73Y128_SLICE_X111Y128_F7BMUX_O),
.O5(CLBLM_L_X72Y128_SLICE_X109Y128_DO5),
.O6(CLBLM_L_X72Y128_SLICE_X109Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33663c3c99cc3c3c)
  ) CLBLM_L_X72Y128_SLICE_X109Y128_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(CLBLL_L_X2Y123_SLICE_X0Y123_CO6),
.I2(CLBLL_R_X73Y128_SLICE_X110Y128_F8MUX_O),
.I3(CLBLM_L_X72Y128_SLICE_X109Y128_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLL_R_X73Y128_SLICE_X111Y128_F7AMUX_O),
.O5(CLBLM_L_X72Y128_SLICE_X109Y128_CO5),
.O6(CLBLM_L_X72Y128_SLICE_X109Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaa00aa)
  ) CLBLM_L_X72Y128_SLICE_X109Y128_BLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y128_SLICE_X109Y128_BO5),
.O6(CLBLM_L_X72Y128_SLICE_X109Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefec2f2ce3e02320)
  ) CLBLM_L_X72Y128_SLICE_X109Y128_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I4(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.O5(CLBLM_L_X72Y128_SLICE_X109Y128_AO5),
.O6(CLBLM_L_X72Y128_SLICE_X109Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y128_SLICE_X109Y128_MUXF7A (
.I0(CLBLM_L_X72Y128_SLICE_X109Y128_BO6),
.I1(CLBLM_L_X72Y128_SLICE_X109Y128_AO6),
.O(CLBLM_L_X72Y128_SLICE_X109Y128_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_DLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X72Y129_SLICE_X108Y129_DO5),
.O6(CLBLM_L_X72Y129_SLICE_X108Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe3ece02f232c20)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_CLUT (
.I0(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I4(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.O5(CLBLM_L_X72Y129_SLICE_X108Y129_CO5),
.O6(CLBLM_L_X72Y129_SLICE_X108Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaf0f0ff00)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_BLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I1(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y129_SLICE_X108Y129_BO5),
.O6(CLBLM_L_X72Y129_SLICE_X108Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haffcaf0ca0fca00c)
  ) CLBLM_L_X72Y129_SLICE_X108Y129_ALUT (
.I0(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.O5(CLBLM_L_X72Y129_SLICE_X108Y129_AO5),
.O6(CLBLM_L_X72Y129_SLICE_X108Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y129_SLICE_X108Y129_MUXF7A (
.I0(CLBLM_L_X72Y129_SLICE_X108Y129_BO6),
.I1(CLBLM_L_X72Y129_SLICE_X108Y129_AO6),
.O(CLBLM_L_X72Y129_SLICE_X108Y129_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y129_SLICE_X108Y129_MUXF7B (
.I0(CLBLM_L_X72Y129_SLICE_X108Y129_DO6),
.I1(CLBLM_L_X72Y129_SLICE_X108Y129_CO6),
.O(CLBLM_L_X72Y129_SLICE_X108Y129_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X72Y129_SLICE_X108Y129_MUXF8 (
.I0(CLBLM_L_X72Y129_SLICE_X108Y129_F7BMUX_O),
.I1(CLBLM_L_X72Y129_SLICE_X108Y129_F7AMUX_O),
.O(CLBLM_L_X72Y129_SLICE_X108Y129_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff00cccc)
  ) CLBLM_L_X72Y129_SLICE_X109Y129_DLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X72Y129_SLICE_X109Y129_DO5),
.O6(CLBLM_L_X72Y129_SLICE_X109Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500e4e4e4e4)
  ) CLBLM_L_X72Y129_SLICE_X109Y129_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I2(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I4(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X72Y129_SLICE_X109Y129_CO5),
.O6(CLBLM_L_X72Y129_SLICE_X109Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbd97351eac86240)
  ) CLBLM_L_X72Y129_SLICE_X109Y129_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I5(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.O5(CLBLM_L_X72Y129_SLICE_X109Y129_BO5),
.O6(CLBLM_L_X72Y129_SLICE_X109Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fa0afa0a)
  ) CLBLM_L_X72Y129_SLICE_X109Y129_ALUT (
.I0(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X72Y129_SLICE_X109Y129_AO5),
.O6(CLBLM_L_X72Y129_SLICE_X109Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y129_SLICE_X109Y129_MUXF7A (
.I0(CLBLM_L_X72Y129_SLICE_X109Y129_BO6),
.I1(CLBLM_L_X72Y129_SLICE_X109Y129_AO6),
.O(CLBLM_L_X72Y129_SLICE_X109Y129_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X72Y129_SLICE_X109Y129_MUXF7B (
.I0(CLBLM_L_X72Y129_SLICE_X109Y129_DO6),
.I1(CLBLM_L_X72Y129_SLICE_X109Y129_CO6),
.O(CLBLM_L_X72Y129_SLICE_X109Y129_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLL_R_X71Y131_SLICE_X107Y131_AO6),
.Q(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb9694da24eb83297)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_DLUT (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I1(CLBLM_L_X72Y128_SLICE_X109Y128_CO6),
.I2(CLBLM_L_X74Y128_SLICE_X112Y128_CO6),
.I3(CLBLL_R_X73Y129_SLICE_X110Y129_CO6),
.I4(CLBLM_L_X72Y128_SLICE_X109Y128_DO6),
.I5(CLBLL_R_X75Y127_SLICE_X114Y127_CO6),
.O5(CLBLM_L_X72Y131_SLICE_X108Y131_DO5),
.O6(CLBLM_L_X72Y131_SLICE_X108Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h21d76e349929a4db)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_CLUT (
.I0(CLBLL_R_X75Y128_SLICE_X115Y128_CO6),
.I1(CLBLM_L_X72Y128_SLICE_X109Y128_CO6),
.I2(CLBLM_L_X74Y128_SLICE_X112Y128_CO6),
.I3(CLBLL_R_X73Y129_SLICE_X110Y129_CO6),
.I4(CLBLM_L_X72Y128_SLICE_X109Y128_DO6),
.I5(CLBLL_R_X75Y127_SLICE_X114Y127_CO6),
.O5(CLBLM_L_X72Y131_SLICE_X108Y131_CO5),
.O6(CLBLM_L_X72Y131_SLICE_X108Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffedffe8004d0048)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(CLBLL_R_X71Y131_SLICE_X107Y131_CQ),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.I4(RIOB33_X105Y169_IOB_X1Y170_I),
.I5(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.O5(CLBLM_L_X72Y131_SLICE_X108Y131_BO5),
.O6(CLBLM_L_X72Y131_SLICE_X108Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a596a)
  ) CLBLM_L_X72Y131_SLICE_X108Y131_ALUT (
.I0(CLBLM_L_X72Y131_SLICE_X108Y131_DO6),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLM_L_X72Y131_SLICE_X108Y131_AQ),
.I3(CLBLM_L_X72Y131_SLICE_X108Y131_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(LIOB33_X0Y79_IOB_X0Y80_I),
.O5(CLBLM_L_X72Y131_SLICE_X108Y131_AO5),
.O6(CLBLM_L_X72Y131_SLICE_X108Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y131_SLICE_X109Y131_DO5),
.O6(CLBLM_L_X72Y131_SLICE_X109Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y131_SLICE_X109Y131_CO5),
.O6(CLBLM_L_X72Y131_SLICE_X109Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y131_SLICE_X109Y131_BO5),
.O6(CLBLM_L_X72Y131_SLICE_X109Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X72Y131_SLICE_X109Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X72Y131_SLICE_X109Y131_AO5),
.O6(CLBLM_L_X72Y131_SLICE_X109Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y115_SLICE_X112Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y115_SLICE_X112Y115_DO5),
.O6(CLBLM_L_X74Y115_SLICE_X112Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y115_SLICE_X112Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y115_SLICE_X112Y115_CO5),
.O6(CLBLM_L_X74Y115_SLICE_X112Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y115_SLICE_X112Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y115_SLICE_X112Y115_BO5),
.O6(CLBLM_L_X74Y115_SLICE_X112Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y115_SLICE_X112Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y115_SLICE_X112Y115_AO5),
.O6(CLBLM_L_X74Y115_SLICE_X112Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfafcfa0c0afc0a0)
  ) CLBLM_L_X74Y115_SLICE_X113Y115_DLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I5(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.O5(CLBLM_L_X74Y115_SLICE_X113Y115_DO5),
.O6(CLBLM_L_X74Y115_SLICE_X113Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef4fea4ae545e040)
  ) CLBLM_L_X74Y115_SLICE_X113Y115_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I5(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.O5(CLBLM_L_X74Y115_SLICE_X113Y115_CO5),
.O6(CLBLM_L_X74Y115_SLICE_X113Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ccaa00f0ccaa)
  ) CLBLM_L_X74Y115_SLICE_X113Y115_BLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.O5(CLBLM_L_X74Y115_SLICE_X113Y115_BO5),
.O6(CLBLM_L_X74Y115_SLICE_X113Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfff0aacc00f0aa)
  ) CLBLM_L_X74Y115_SLICE_X113Y115_ALUT (
.I0(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.O5(CLBLM_L_X74Y115_SLICE_X113Y115_AO5),
.O6(CLBLM_L_X74Y115_SLICE_X113Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y115_SLICE_X113Y115_MUXF7A (
.I0(CLBLM_L_X74Y115_SLICE_X113Y115_BO6),
.I1(CLBLM_L_X74Y115_SLICE_X113Y115_AO6),
.O(CLBLM_L_X74Y115_SLICE_X113Y115_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y115_SLICE_X113Y115_MUXF7B (
.I0(CLBLM_L_X74Y115_SLICE_X113Y115_DO6),
.I1(CLBLM_L_X74Y115_SLICE_X113Y115_CO6),
.O(CLBLM_L_X74Y115_SLICE_X113Y115_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y115_SLICE_X113Y115_MUXF8 (
.I0(CLBLM_L_X74Y115_SLICE_X113Y115_F7BMUX_O),
.I1(CLBLM_L_X74Y115_SLICE_X113Y115_F7AMUX_O),
.O(CLBLM_L_X74Y115_SLICE_X113Y115_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dd88dd88)
  ) CLBLM_L_X74Y116_SLICE_X112Y116_DLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I4(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X74Y116_SLICE_X112Y116_DO5),
.O6(CLBLM_L_X74Y116_SLICE_X112Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaef4a45e0e5404)
  ) CLBLM_L_X74Y116_SLICE_X112Y116_CLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I5(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.O5(CLBLM_L_X74Y116_SLICE_X112Y116_CO5),
.O6(CLBLM_L_X74Y116_SLICE_X112Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe5ef454ae0ea404)
  ) CLBLM_L_X74Y116_SLICE_X112Y116_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.O5(CLBLM_L_X74Y116_SLICE_X112Y116_BO5),
.O6(CLBLM_L_X74Y116_SLICE_X112Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cfcfafa0c0c0)
  ) CLBLM_L_X74Y116_SLICE_X112Y116_ALUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.O5(CLBLM_L_X74Y116_SLICE_X112Y116_AO5),
.O6(CLBLM_L_X74Y116_SLICE_X112Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y116_SLICE_X112Y116_MUXF7A (
.I0(CLBLM_L_X74Y116_SLICE_X112Y116_BO6),
.I1(CLBLM_L_X74Y116_SLICE_X112Y116_AO6),
.O(CLBLM_L_X74Y116_SLICE_X112Y116_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y116_SLICE_X112Y116_MUXF7B (
.I0(CLBLM_L_X74Y116_SLICE_X112Y116_DO6),
.I1(CLBLM_L_X74Y116_SLICE_X112Y116_CO6),
.O(CLBLM_L_X74Y116_SLICE_X112Y116_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y116_SLICE_X112Y116_MUXF8 (
.I0(CLBLM_L_X74Y116_SLICE_X112Y116_F7BMUX_O),
.I1(CLBLM_L_X74Y116_SLICE_X112Y116_F7AMUX_O),
.O(CLBLM_L_X74Y116_SLICE_X112Y116_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y116_SLICE_X113Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y116_SLICE_X113Y116_DO5),
.O6(CLBLM_L_X74Y116_SLICE_X113Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f4b3c7887c3b4f0)
  ) CLBLM_L_X74Y116_SLICE_X113Y116_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(CLBLM_L_X70Y121_SLICE_X104Y121_DO6),
.I3(CLBLM_L_X74Y116_SLICE_X113Y116_F7AMUX_O),
.I4(CLBLM_L_X74Y115_SLICE_X113Y115_F8MUX_O),
.I5(CLBLL_R_X75Y116_SLICE_X115Y116_F7AMUX_O),
.O5(CLBLM_L_X74Y116_SLICE_X113Y116_CO5),
.O6(CLBLM_L_X74Y116_SLICE_X113Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfa0a0c0cfa0a)
  ) CLBLM_L_X74Y116_SLICE_X113Y116_BLUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I1(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLM_L_X74Y116_SLICE_X113Y116_BO5),
.O6(CLBLM_L_X74Y116_SLICE_X113Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd75b931ec64a820)
  ) CLBLM_L_X74Y116_SLICE_X113Y116_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I4(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.O5(CLBLM_L_X74Y116_SLICE_X113Y116_AO5),
.O6(CLBLM_L_X74Y116_SLICE_X113Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y116_SLICE_X113Y116_MUXF7A (
.I0(CLBLM_L_X74Y116_SLICE_X113Y116_BO6),
.I1(CLBLM_L_X74Y116_SLICE_X113Y116_AO6),
.O(CLBLM_L_X74Y116_SLICE_X113Y116_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcce2e23300e2e2)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_DLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I3(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.O5(CLBLM_L_X74Y117_SLICE_X112Y117_DO5),
.O6(CLBLM_L_X74Y117_SLICE_X112Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeef5a04444f5a0)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.O5(CLBLM_L_X74Y117_SLICE_X112Y117_CO5),
.O6(CLBLM_L_X74Y117_SLICE_X112Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbea7362d9c85140)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I4(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.O5(CLBLM_L_X74Y117_SLICE_X112Y117_BO5),
.O6(CLBLM_L_X74Y117_SLICE_X112Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaae4e45500e4e4)
  ) CLBLM_L_X74Y117_SLICE_X112Y117_ALUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I3(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.O5(CLBLM_L_X74Y117_SLICE_X112Y117_AO5),
.O6(CLBLM_L_X74Y117_SLICE_X112Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y117_SLICE_X112Y117_MUXF7A (
.I0(CLBLM_L_X74Y117_SLICE_X112Y117_BO6),
.I1(CLBLM_L_X74Y117_SLICE_X112Y117_AO6),
.O(CLBLM_L_X74Y117_SLICE_X112Y117_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y117_SLICE_X112Y117_MUXF7B (
.I0(CLBLM_L_X74Y117_SLICE_X112Y117_DO6),
.I1(CLBLM_L_X74Y117_SLICE_X112Y117_CO6),
.O(CLBLM_L_X74Y117_SLICE_X112Y117_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y117_SLICE_X112Y117_MUXF8 (
.I0(CLBLM_L_X74Y117_SLICE_X112Y117_F7BMUX_O),
.I1(CLBLM_L_X74Y117_SLICE_X112Y117_F7AMUX_O),
.O(CLBLM_L_X74Y117_SLICE_X112Y117_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2075df8a2a7fd580)
  ) CLBLM_L_X74Y117_SLICE_X113Y117_DLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLM_L_X74Y118_SLICE_X113Y118_F7AMUX_O),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(CLBLL_R_X75Y117_SLICE_X115Y117_F8MUX_O),
.I4(CLBLM_L_X70Y121_SLICE_X104Y121_DO6),
.I5(CLBLL_R_X75Y117_SLICE_X114Y117_F7BMUX_O),
.O5(CLBLM_L_X74Y117_SLICE_X113Y117_DO5),
.O6(CLBLM_L_X74Y117_SLICE_X113Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3636369c9c9c369c)
  ) CLBLM_L_X74Y117_SLICE_X113Y117_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y82_I),
.I1(CLBLL_R_X71Y131_SLICE_X107Y131_AO6),
.I2(CLBLM_L_X74Y117_SLICE_X112Y117_F8MUX_O),
.I3(CLBLM_L_X74Y117_SLICE_X113Y117_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_R_X75Y117_SLICE_X114Y117_F7AMUX_O),
.O5(CLBLM_L_X74Y117_SLICE_X113Y117_CO5),
.O6(CLBLM_L_X74Y117_SLICE_X113Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cafaffc0ca0a0)
  ) CLBLM_L_X74Y117_SLICE_X113Y117_BLUT (
.I0(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.O5(CLBLM_L_X74Y117_SLICE_X113Y117_BO5),
.O6(CLBLM_L_X74Y117_SLICE_X113Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfadd5088fa8850)
  ) CLBLM_L_X74Y117_SLICE_X113Y117_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.O5(CLBLM_L_X74Y117_SLICE_X113Y117_AO5),
.O6(CLBLM_L_X74Y117_SLICE_X113Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y117_SLICE_X113Y117_MUXF7A (
.I0(CLBLM_L_X74Y117_SLICE_X113Y117_BO6),
.I1(CLBLM_L_X74Y117_SLICE_X113Y117_AO6),
.O(CLBLM_L_X74Y117_SLICE_X113Y117_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X112Y118_DO5),
.O6(CLBLM_L_X74Y118_SLICE_X112Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X112Y118_CO5),
.O6(CLBLM_L_X74Y118_SLICE_X112Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X112Y118_BO5),
.O6(CLBLM_L_X74Y118_SLICE_X112Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X112Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X112Y118_AO5),
.O6(CLBLM_L_X74Y118_SLICE_X112Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X113Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X113Y118_DO5),
.O6(CLBLM_L_X74Y118_SLICE_X113Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y118_SLICE_X113Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y118_SLICE_X113Y118_CO5),
.O6(CLBLM_L_X74Y118_SLICE_X113Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef4fea4ae545e040)
  ) CLBLM_L_X74Y118_SLICE_X113Y118_BLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I4(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.O5(CLBLM_L_X74Y118_SLICE_X113Y118_BO5),
.O6(CLBLM_L_X74Y118_SLICE_X113Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfd58f85dad08a80)
  ) CLBLM_L_X74Y118_SLICE_X113Y118_ALUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I5(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.O5(CLBLM_L_X74Y118_SLICE_X113Y118_AO5),
.O6(CLBLM_L_X74Y118_SLICE_X113Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y118_SLICE_X113Y118_MUXF7A (
.I0(CLBLM_L_X74Y118_SLICE_X113Y118_BO6),
.I1(CLBLM_L_X74Y118_SLICE_X113Y118_AO6),
.O(CLBLM_L_X74Y118_SLICE_X113Y118_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaee445050ee44)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_DLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.O5(CLBLM_L_X74Y119_SLICE_X112Y119_DO5),
.O6(CLBLM_L_X74Y119_SLICE_X112Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe455e4aae400e4)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.O5(CLBLM_L_X74Y119_SLICE_X112Y119_CO5),
.O6(CLBLM_L_X74Y119_SLICE_X112Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacff0facacf000)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_BLUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.O5(CLBLM_L_X74Y119_SLICE_X112Y119_BO5),
.O6(CLBLM_L_X74Y119_SLICE_X112Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0fafacfc00a0a)
  ) CLBLM_L_X74Y119_SLICE_X112Y119_ALUT (
.I0(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.O5(CLBLM_L_X74Y119_SLICE_X112Y119_AO5),
.O6(CLBLM_L_X74Y119_SLICE_X112Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y119_SLICE_X112Y119_MUXF7A (
.I0(CLBLM_L_X74Y119_SLICE_X112Y119_BO6),
.I1(CLBLM_L_X74Y119_SLICE_X112Y119_AO6),
.O(CLBLM_L_X74Y119_SLICE_X112Y119_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y119_SLICE_X112Y119_MUXF7B (
.I0(CLBLM_L_X74Y119_SLICE_X112Y119_DO6),
.I1(CLBLM_L_X74Y119_SLICE_X112Y119_CO6),
.O(CLBLM_L_X74Y119_SLICE_X112Y119_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y119_SLICE_X112Y119_MUXF8 (
.I0(CLBLM_L_X74Y119_SLICE_X112Y119_F7BMUX_O),
.I1(CLBLM_L_X74Y119_SLICE_X112Y119_F7AMUX_O),
.O(CLBLM_L_X74Y119_SLICE_X112Y119_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacaff0fcacaf000)
  ) CLBLM_L_X74Y119_SLICE_X113Y119_DLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLM_L_X74Y119_SLICE_X113Y119_DO5),
.O6(CLBLM_L_X74Y119_SLICE_X113Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf8fbc8cb383b080)
  ) CLBLM_L_X74Y119_SLICE_X113Y119_CLUT (
.I0(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I1(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.O5(CLBLM_L_X74Y119_SLICE_X113Y119_CO5),
.O6(CLBLM_L_X74Y119_SLICE_X113Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaaaff00)
  ) CLBLM_L_X74Y119_SLICE_X113Y119_BLUT (
.I0(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLM_L_X74Y119_SLICE_X113Y119_BO5),
.O6(CLBLM_L_X74Y119_SLICE_X113Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfafc0afcfa0c0a0)
  ) CLBLM_L_X74Y119_SLICE_X113Y119_ALUT (
.I0(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.O5(CLBLM_L_X74Y119_SLICE_X113Y119_AO5),
.O6(CLBLM_L_X74Y119_SLICE_X113Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y119_SLICE_X113Y119_MUXF7A (
.I0(CLBLM_L_X74Y119_SLICE_X113Y119_BO6),
.I1(CLBLM_L_X74Y119_SLICE_X113Y119_AO6),
.O(CLBLM_L_X74Y119_SLICE_X113Y119_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y119_SLICE_X113Y119_MUXF7B (
.I0(CLBLM_L_X74Y119_SLICE_X113Y119_DO6),
.I1(CLBLM_L_X74Y119_SLICE_X113Y119_CO6),
.O(CLBLM_L_X74Y119_SLICE_X113Y119_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccf0ffaaccf000)
  ) CLBLM_L_X74Y120_SLICE_X112Y120_DLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.I2(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.O5(CLBLM_L_X74Y120_SLICE_X112Y120_DO5),
.O6(CLBLM_L_X74Y120_SLICE_X112Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4ffe4aae455e400)
  ) CLBLM_L_X74Y120_SLICE_X112Y120_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.O5(CLBLM_L_X74Y120_SLICE_X112Y120_CO5),
.O6(CLBLM_L_X74Y120_SLICE_X112Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44f5f5a0a0)
  ) CLBLM_L_X74Y120_SLICE_X112Y120_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLM_L_X74Y120_SLICE_X112Y120_BO5),
.O6(CLBLM_L_X74Y120_SLICE_X112Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5dd88a0a0dd88)
  ) CLBLM_L_X74Y120_SLICE_X112Y120_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I2(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I3(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.O5(CLBLM_L_X74Y120_SLICE_X112Y120_AO5),
.O6(CLBLM_L_X74Y120_SLICE_X112Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y120_SLICE_X112Y120_MUXF7A (
.I0(CLBLM_L_X74Y120_SLICE_X112Y120_BO6),
.I1(CLBLM_L_X74Y120_SLICE_X112Y120_AO6),
.O(CLBLM_L_X74Y120_SLICE_X112Y120_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y120_SLICE_X112Y120_MUXF7B (
.I0(CLBLM_L_X74Y120_SLICE_X112Y120_DO6),
.I1(CLBLM_L_X74Y120_SLICE_X112Y120_CO6),
.O(CLBLM_L_X74Y120_SLICE_X112Y120_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y120_SLICE_X112Y120_MUXF8 (
.I0(CLBLM_L_X74Y120_SLICE_X112Y120_F7BMUX_O),
.I1(CLBLM_L_X74Y120_SLICE_X112Y120_F7AMUX_O),
.O(CLBLM_L_X74Y120_SLICE_X112Y120_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y120_SLICE_X113Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y120_SLICE_X113Y120_DO5),
.O6(CLBLM_L_X74Y120_SLICE_X113Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y120_SLICE_X113Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y120_SLICE_X113Y120_CO5),
.O6(CLBLM_L_X74Y120_SLICE_X113Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y120_SLICE_X113Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y120_SLICE_X113Y120_BO5),
.O6(CLBLM_L_X74Y120_SLICE_X113Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c3f5555f3c0aaaa)
  ) CLBLM_L_X74Y120_SLICE_X113Y120_ALUT (
.I0(CLBLM_L_X74Y121_SLICE_X113Y121_F8MUX_O),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(CLBLM_L_X74Y119_SLICE_X113Y119_F7BMUX_O),
.I3(CLBLM_L_X74Y119_SLICE_X113Y119_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.O5(CLBLM_L_X74Y120_SLICE_X113Y120_AO5),
.O6(CLBLM_L_X74Y120_SLICE_X113Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfa88fadd508850)
  ) CLBLM_L_X74Y121_SLICE_X112Y121_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.I3(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I4(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.O5(CLBLM_L_X74Y121_SLICE_X112Y121_DO5),
.O6(CLBLM_L_X74Y121_SLICE_X112Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30eeeefc302222)
  ) CLBLM_L_X74Y121_SLICE_X112Y121_CLUT (
.I0(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I4(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.O5(CLBLM_L_X74Y121_SLICE_X112Y121_CO5),
.O6(CLBLM_L_X74Y121_SLICE_X112Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4ff55e4e4aa00)
  ) CLBLM_L_X74Y121_SLICE_X112Y121_BLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I3(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.O5(CLBLM_L_X74Y121_SLICE_X112Y121_BO5),
.O6(CLBLM_L_X74Y121_SLICE_X112Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd5df858ad0da808)
  ) CLBLM_L_X74Y121_SLICE_X112Y121_ALUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.O5(CLBLM_L_X74Y121_SLICE_X112Y121_AO5),
.O6(CLBLM_L_X74Y121_SLICE_X112Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y121_SLICE_X112Y121_MUXF7A (
.I0(CLBLM_L_X74Y121_SLICE_X112Y121_BO6),
.I1(CLBLM_L_X74Y121_SLICE_X112Y121_AO6),
.O(CLBLM_L_X74Y121_SLICE_X112Y121_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y121_SLICE_X112Y121_MUXF7B (
.I0(CLBLM_L_X74Y121_SLICE_X112Y121_DO6),
.I1(CLBLM_L_X74Y121_SLICE_X112Y121_CO6),
.O(CLBLM_L_X74Y121_SLICE_X112Y121_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y121_SLICE_X112Y121_MUXF8 (
.I0(CLBLM_L_X74Y121_SLICE_X112Y121_F7BMUX_O),
.I1(CLBLM_L_X74Y121_SLICE_X112Y121_F7AMUX_O),
.O(CLBLM_L_X74Y121_SLICE_X112Y121_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcaffca00caf0ca0)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_DLUT (
.I0(CLBLL_R_X77Y113_SLICE_X118Y113_CO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_CO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I5(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.O5(CLBLM_L_X74Y121_SLICE_X113Y121_DO5),
.O6(CLBLM_L_X74Y121_SLICE_X113Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffac0facf0ac00ac)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_CLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_BO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_BO6),
.I2(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_BO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_BO6),
.O5(CLBLM_L_X74Y121_SLICE_X113Y121_CO5),
.O6(CLBLM_L_X74Y121_SLICE_X113Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdecb9a875643120)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_BLUT (
.I0(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y126_SLICE_X120Y126_AO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_BO6),
.I4(CLBLM_L_X78Y121_SLICE_X120Y121_AO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_BO6),
.O5(CLBLM_L_X74Y121_SLICE_X113Y121_BO5),
.O6(CLBLM_L_X74Y121_SLICE_X113Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaf0ccf0cc)
  ) CLBLM_L_X74Y121_SLICE_X113Y121_ALUT (
.I0(CLBLL_R_X77Y115_SLICE_X118Y115_AO6),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I2(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_DO6),
.I5(CLBLL_R_X73Y119_SLICE_X111Y119_DO6),
.O5(CLBLM_L_X74Y121_SLICE_X113Y121_AO5),
.O6(CLBLM_L_X74Y121_SLICE_X113Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y121_SLICE_X113Y121_MUXF7A (
.I0(CLBLM_L_X74Y121_SLICE_X113Y121_BO6),
.I1(CLBLM_L_X74Y121_SLICE_X113Y121_AO6),
.O(CLBLM_L_X74Y121_SLICE_X113Y121_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y121_SLICE_X113Y121_MUXF7B (
.I0(CLBLM_L_X74Y121_SLICE_X113Y121_DO6),
.I1(CLBLM_L_X74Y121_SLICE_X113Y121_CO6),
.O(CLBLM_L_X74Y121_SLICE_X113Y121_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y121_SLICE_X113Y121_MUXF8 (
.I0(CLBLM_L_X74Y121_SLICE_X113Y121_F7BMUX_O),
.I1(CLBLM_L_X74Y121_SLICE_X113Y121_F7AMUX_O),
.O(CLBLM_L_X74Y121_SLICE_X113Y121_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y123_SLICE_X112Y123_DO5),
.O6(CLBLM_L_X74Y123_SLICE_X112Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc3c3c66663c3c)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_CLUT (
.I0(CLBLM_L_X74Y124_SLICE_X113Y124_F7BMUX_O),
.I1(CLBLL_R_X71Y128_SLICE_X106Y128_CO6),
.I2(CLBLM_L_X74Y123_SLICE_X113Y123_F8MUX_O),
.I3(CLBLM_L_X74Y125_SLICE_X112Y125_F7AMUX_O),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_L_X74Y123_SLICE_X112Y123_CO5),
.O6(CLBLM_L_X74Y123_SLICE_X112Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8ffaad8d85500)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I2(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.O5(CLBLM_L_X74Y123_SLICE_X112Y123_BO5),
.O6(CLBLM_L_X74Y123_SLICE_X112Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5eea0eef544a044)
  ) CLBLM_L_X74Y123_SLICE_X112Y123_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.O5(CLBLM_L_X74Y123_SLICE_X112Y123_AO5),
.O6(CLBLM_L_X74Y123_SLICE_X112Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y123_SLICE_X112Y123_MUXF7A (
.I0(CLBLM_L_X74Y123_SLICE_X112Y123_BO6),
.I1(CLBLM_L_X74Y123_SLICE_X112Y123_AO6),
.O(CLBLM_L_X74Y123_SLICE_X112Y123_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0fff000)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_DLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I1(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X74Y123_SLICE_X113Y123_DO5),
.O6(CLBLM_L_X74Y123_SLICE_X113Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cafafa0a0)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_CLUT (
.I0(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I1(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X74Y123_SLICE_X113Y123_CO5),
.O6(CLBLM_L_X74Y123_SLICE_X113Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd8aad855d800d8)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I2(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.O5(CLBLM_L_X74Y123_SLICE_X113Y123_BO5),
.O6(CLBLM_L_X74Y123_SLICE_X113Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe76ba32dc549810)
  ) CLBLM_L_X74Y123_SLICE_X113Y123_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.O5(CLBLM_L_X74Y123_SLICE_X113Y123_AO5),
.O6(CLBLM_L_X74Y123_SLICE_X113Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y123_SLICE_X113Y123_MUXF7A (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_BO6),
.I1(CLBLM_L_X74Y123_SLICE_X113Y123_AO6),
.O(CLBLM_L_X74Y123_SLICE_X113Y123_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y123_SLICE_X113Y123_MUXF7B (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_DO6),
.I1(CLBLM_L_X74Y123_SLICE_X113Y123_CO6),
.O(CLBLM_L_X74Y123_SLICE_X113Y123_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y123_SLICE_X113Y123_MUXF8 (
.I0(CLBLM_L_X74Y123_SLICE_X113Y123_F7BMUX_O),
.I1(CLBLM_L_X74Y123_SLICE_X113Y123_F7AMUX_O),
.O(CLBLM_L_X74Y123_SLICE_X113Y123_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccf0ffaaccf000)
  ) CLBLM_L_X74Y124_SLICE_X112Y124_DLUT (
.I0(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I2(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.O5(CLBLM_L_X74Y124_SLICE_X112Y124_DO5),
.O6(CLBLM_L_X74Y124_SLICE_X112Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0fff000)
  ) CLBLM_L_X74Y124_SLICE_X112Y124_CLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X74Y124_SLICE_X112Y124_CO5),
.O6(CLBLM_L_X74Y124_SLICE_X112Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0fafacfc00a0a)
  ) CLBLM_L_X74Y124_SLICE_X112Y124_BLUT (
.I0(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.O5(CLBLM_L_X74Y124_SLICE_X112Y124_BO5),
.O6(CLBLM_L_X74Y124_SLICE_X112Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3eef322c0eec022)
  ) CLBLM_L_X74Y124_SLICE_X112Y124_ALUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.O5(CLBLM_L_X74Y124_SLICE_X112Y124_AO5),
.O6(CLBLM_L_X74Y124_SLICE_X112Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y124_SLICE_X112Y124_MUXF7A (
.I0(CLBLM_L_X74Y124_SLICE_X112Y124_BO6),
.I1(CLBLM_L_X74Y124_SLICE_X112Y124_AO6),
.O(CLBLM_L_X74Y124_SLICE_X112Y124_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y124_SLICE_X112Y124_MUXF7B (
.I0(CLBLM_L_X74Y124_SLICE_X112Y124_DO6),
.I1(CLBLM_L_X74Y124_SLICE_X112Y124_CO6),
.O(CLBLM_L_X74Y124_SLICE_X112Y124_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y124_SLICE_X112Y124_MUXF8 (
.I0(CLBLM_L_X74Y124_SLICE_X112Y124_F7BMUX_O),
.I1(CLBLM_L_X74Y124_SLICE_X112Y124_F7AMUX_O),
.O(CLBLM_L_X74Y124_SLICE_X112Y124_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf8ada85d580d08)
  ) CLBLM_L_X74Y124_SLICE_X113Y124_DLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.O5(CLBLM_L_X74Y124_SLICE_X113Y124_DO5),
.O6(CLBLM_L_X74Y124_SLICE_X113Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haffca0fcaf0ca00c)
  ) CLBLM_L_X74Y124_SLICE_X113Y124_CLUT (
.I0(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I5(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.O5(CLBLM_L_X74Y124_SLICE_X113Y124_CO5),
.O6(CLBLM_L_X74Y124_SLICE_X113Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaa00aa)
  ) CLBLM_L_X74Y124_SLICE_X113Y124_BLUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I2(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X74Y124_SLICE_X113Y124_BO5),
.O6(CLBLM_L_X74Y124_SLICE_X113Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbd97351eac86240)
  ) CLBLM_L_X74Y124_SLICE_X113Y124_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.O5(CLBLM_L_X74Y124_SLICE_X113Y124_AO5),
.O6(CLBLM_L_X74Y124_SLICE_X113Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y124_SLICE_X113Y124_MUXF7A (
.I0(CLBLM_L_X74Y124_SLICE_X113Y124_BO6),
.I1(CLBLM_L_X74Y124_SLICE_X113Y124_AO6),
.O(CLBLM_L_X74Y124_SLICE_X113Y124_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y124_SLICE_X113Y124_MUXF7B (
.I0(CLBLM_L_X74Y124_SLICE_X113Y124_DO6),
.I1(CLBLM_L_X74Y124_SLICE_X113Y124_CO6),
.O(CLBLM_L_X74Y124_SLICE_X113Y124_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2070df8f2f7fd080)
  ) CLBLM_L_X74Y125_SLICE_X112Y125_DLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(CLBLM_L_X74Y125_SLICE_X113Y125_F7BMUX_O),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(CLBLM_L_X74Y124_SLICE_X113Y124_F7AMUX_O),
.I4(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.I5(CLBLL_R_X73Y125_SLICE_X111Y125_F8MUX_O),
.O5(CLBLM_L_X74Y125_SLICE_X112Y125_DO5),
.O6(CLBLM_L_X74Y125_SLICE_X112Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05f5fa0a3535caca)
  ) CLBLM_L_X74Y125_SLICE_X112Y125_CLUT (
.I0(CLBLM_L_X74Y126_SLICE_X112Y126_F8MUX_O),
.I1(CLBLM_L_X74Y125_SLICE_X113Y125_F7AMUX_O),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(CLBLL_R_X73Y126_SLICE_X111Y126_F7AMUX_O),
.I4(CLBLM_R_X59Y117_SLICE_X88Y117_AO6),
.I5(LIOB33_X0Y81_IOB_X0Y81_I),
.O5(CLBLM_L_X74Y125_SLICE_X112Y125_CO5),
.O6(CLBLM_L_X74Y125_SLICE_X112Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef2fe323ec2ce020)
  ) CLBLM_L_X74Y125_SLICE_X112Y125_BLUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I4(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.O5(CLBLM_L_X74Y125_SLICE_X112Y125_BO5),
.O6(CLBLM_L_X74Y125_SLICE_X112Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccf0ffaaccf000)
  ) CLBLM_L_X74Y125_SLICE_X112Y125_ALUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.O5(CLBLM_L_X74Y125_SLICE_X112Y125_AO5),
.O6(CLBLM_L_X74Y125_SLICE_X112Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y125_SLICE_X112Y125_MUXF7A (
.I0(CLBLM_L_X74Y125_SLICE_X112Y125_BO6),
.I1(CLBLM_L_X74Y125_SLICE_X112Y125_AO6),
.O(CLBLM_L_X74Y125_SLICE_X112Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0cfcfafa0c0c0)
  ) CLBLM_L_X74Y125_SLICE_X113Y125_DLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I4(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.O5(CLBLM_L_X74Y125_SLICE_X113Y125_DO5),
.O6(CLBLM_L_X74Y125_SLICE_X113Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcaffca00caf0ca0)
  ) CLBLM_L_X74Y125_SLICE_X113Y125_CLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I5(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.O5(CLBLM_L_X74Y125_SLICE_X113Y125_CO5),
.O6(CLBLM_L_X74Y125_SLICE_X113Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44f5f5a0a0)
  ) CLBLM_L_X74Y125_SLICE_X113Y125_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I2(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I3(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X74Y125_SLICE_X113Y125_BO5),
.O6(CLBLM_L_X74Y125_SLICE_X113Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0afc0cfc0c)
  ) CLBLM_L_X74Y125_SLICE_X113Y125_ALUT (
.I0(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I4(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X74Y125_SLICE_X113Y125_AO5),
.O6(CLBLM_L_X74Y125_SLICE_X113Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y125_SLICE_X113Y125_MUXF7A (
.I0(CLBLM_L_X74Y125_SLICE_X113Y125_BO6),
.I1(CLBLM_L_X74Y125_SLICE_X113Y125_AO6),
.O(CLBLM_L_X74Y125_SLICE_X113Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y125_SLICE_X113Y125_MUXF7B (
.I0(CLBLM_L_X74Y125_SLICE_X113Y125_DO6),
.I1(CLBLM_L_X74Y125_SLICE_X113Y125_CO6),
.O(CLBLM_L_X74Y125_SLICE_X113Y125_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccffcc00)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_DLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X74Y126_SLICE_X112Y126_DO5),
.O6(CLBLM_L_X74Y126_SLICE_X112Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88f3f3c0c0)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_CLUT (
.I0(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I3(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X74Y126_SLICE_X112Y126_CO5),
.O6(CLBLM_L_X74Y126_SLICE_X112Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccaaf0aaf0)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_BLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I2(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X74Y126_SLICE_X112Y126_BO5),
.O6(CLBLM_L_X74Y126_SLICE_X112Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaaffaa00)
  ) CLBLM_L_X74Y126_SLICE_X112Y126_ALUT (
.I0(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X74Y126_SLICE_X112Y126_AO5),
.O6(CLBLM_L_X74Y126_SLICE_X112Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y126_SLICE_X112Y126_MUXF7A (
.I0(CLBLM_L_X74Y126_SLICE_X112Y126_BO6),
.I1(CLBLM_L_X74Y126_SLICE_X112Y126_AO6),
.O(CLBLM_L_X74Y126_SLICE_X112Y126_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y126_SLICE_X112Y126_MUXF7B (
.I0(CLBLM_L_X74Y126_SLICE_X112Y126_DO6),
.I1(CLBLM_L_X74Y126_SLICE_X112Y126_CO6),
.O(CLBLM_L_X74Y126_SLICE_X112Y126_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y126_SLICE_X112Y126_MUXF8 (
.I0(CLBLM_L_X74Y126_SLICE_X112Y126_F7BMUX_O),
.I1(CLBLM_L_X74Y126_SLICE_X112Y126_F7AMUX_O),
.O(CLBLM_L_X74Y126_SLICE_X112Y126_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y126_SLICE_X113Y126_DO5),
.O6(CLBLM_L_X74Y126_SLICE_X113Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y126_SLICE_X113Y126_CO5),
.O6(CLBLM_L_X74Y126_SLICE_X113Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y126_SLICE_X113Y126_BO5),
.O6(CLBLM_L_X74Y126_SLICE_X113Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y126_SLICE_X113Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y126_SLICE_X113Y126_AO5),
.O6(CLBLM_L_X74Y126_SLICE_X113Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dd88dd88)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I2(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I4(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X74Y127_SLICE_X112Y127_DO5),
.O6(CLBLM_L_X74Y127_SLICE_X112Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ffaa5500)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X74Y127_SLICE_X112Y127_CO5),
.O6(CLBLM_L_X74Y127_SLICE_X112Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaffc0ca0a0fc0c)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_BLUT (
.I0(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.O5(CLBLM_L_X74Y127_SLICE_X112Y127_BO5),
.O6(CLBLM_L_X74Y127_SLICE_X112Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefec2f2ce3e02320)
  ) CLBLM_L_X74Y127_SLICE_X112Y127_ALUT (
.I0(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.O5(CLBLM_L_X74Y127_SLICE_X112Y127_AO5),
.O6(CLBLM_L_X74Y127_SLICE_X112Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y127_SLICE_X112Y127_MUXF7A (
.I0(CLBLM_L_X74Y127_SLICE_X112Y127_BO6),
.I1(CLBLM_L_X74Y127_SLICE_X112Y127_AO6),
.O(CLBLM_L_X74Y127_SLICE_X112Y127_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y127_SLICE_X112Y127_MUXF7B (
.I0(CLBLM_L_X74Y127_SLICE_X112Y127_DO6),
.I1(CLBLM_L_X74Y127_SLICE_X112Y127_CO6),
.O(CLBLM_L_X74Y127_SLICE_X112Y127_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y127_SLICE_X113Y127_DO5),
.O6(CLBLM_L_X74Y127_SLICE_X113Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y127_SLICE_X113Y127_CO5),
.O6(CLBLM_L_X74Y127_SLICE_X113Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22f3f3ee22c0c0)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_BLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.O5(CLBLM_L_X74Y127_SLICE_X113Y127_BO5),
.O6(CLBLM_L_X74Y127_SLICE_X113Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88f5f5dd88a0a0)
  ) CLBLM_L_X74Y127_SLICE_X113Y127_ALUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I2(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I3(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.O5(CLBLM_L_X74Y127_SLICE_X113Y127_AO5),
.O6(CLBLM_L_X74Y127_SLICE_X113Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y127_SLICE_X113Y127_MUXF7A (
.I0(CLBLM_L_X74Y127_SLICE_X113Y127_BO6),
.I1(CLBLM_L_X74Y127_SLICE_X113Y127_AO6),
.O(CLBLM_L_X74Y127_SLICE_X113Y127_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y128_SLICE_X112Y128_DO5),
.O6(CLBLM_L_X74Y128_SLICE_X112Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h339966cc3c3c3c3c)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_CLUT (
.I0(LIOB33_X0Y81_IOB_X0Y81_I),
.I1(CLBLM_L_X70Y128_SLICE_X105Y128_CO6),
.I2(CLBLL_R_X75Y128_SLICE_X114Y128_F8MUX_O),
.I3(CLBLM_L_X74Y128_SLICE_X112Y128_F7AMUX_O),
.I4(CLBLM_L_X74Y127_SLICE_X112Y127_F7BMUX_O),
.I5(LIOB33_X0Y81_IOB_X0Y82_I),
.O5(CLBLM_L_X74Y128_SLICE_X112Y128_CO5),
.O6(CLBLM_L_X74Y128_SLICE_X112Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88fcfcbb883030)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_BLUT (
.I0(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.O5(CLBLM_L_X74Y128_SLICE_X112Y128_BO5),
.O6(CLBLM_L_X74Y128_SLICE_X112Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_L_X74Y128_SLICE_X112Y128_ALUT (
.I0(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I2(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X74Y128_SLICE_X112Y128_AO5),
.O6(CLBLM_L_X74Y128_SLICE_X112Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y128_SLICE_X112Y128_MUXF7A (
.I0(CLBLM_L_X74Y128_SLICE_X112Y128_BO6),
.I1(CLBLM_L_X74Y128_SLICE_X112Y128_AO6),
.O(CLBLM_L_X74Y128_SLICE_X112Y128_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLM_L_X74Y128_SLICE_X113Y128_DLUT (
.I0(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I1(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I2(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I3(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X74Y128_SLICE_X113Y128_DO5),
.O6(CLBLM_L_X74Y128_SLICE_X113Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050dd88dd88)
  ) CLBLM_L_X74Y128_SLICE_X113Y128_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.I4(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I5(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.O5(CLBLM_L_X74Y128_SLICE_X113Y128_CO5),
.O6(CLBLM_L_X74Y128_SLICE_X113Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefe54f45eae04a40)
  ) CLBLM_L_X74Y128_SLICE_X113Y128_BLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.O5(CLBLM_L_X74Y128_SLICE_X113Y128_BO5),
.O6(CLBLM_L_X74Y128_SLICE_X113Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLM_L_X74Y128_SLICE_X113Y128_ALUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X74Y128_SLICE_X113Y128_AO5),
.O6(CLBLM_L_X74Y128_SLICE_X113Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y128_SLICE_X113Y128_MUXF7A (
.I0(CLBLM_L_X74Y128_SLICE_X113Y128_BO6),
.I1(CLBLM_L_X74Y128_SLICE_X113Y128_AO6),
.O(CLBLM_L_X74Y128_SLICE_X113Y128_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y128_SLICE_X113Y128_MUXF7B (
.I0(CLBLM_L_X74Y128_SLICE_X113Y128_DO6),
.I1(CLBLM_L_X74Y128_SLICE_X113Y128_CO6),
.O(CLBLM_L_X74Y128_SLICE_X113Y128_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X74Y128_SLICE_X113Y128_MUXF8 (
.I0(CLBLM_L_X74Y128_SLICE_X113Y128_F7BMUX_O),
.I1(CLBLM_L_X74Y128_SLICE_X113Y128_F7AMUX_O),
.O(CLBLM_L_X74Y128_SLICE_X113Y128_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X112Y129_DO5),
.O6(CLBLM_L_X74Y129_SLICE_X112Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X112Y129_CO5),
.O6(CLBLM_L_X74Y129_SLICE_X112Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaf0f0cccc)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_BLUT (
.I0(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I2(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.I3(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I4(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X74Y129_SLICE_X112Y129_BO5),
.O6(CLBLM_L_X74Y129_SLICE_X112Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444fa50fa50)
  ) CLBLM_L_X74Y129_SLICE_X112Y129_ALUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I2(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I3(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I4(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X74Y129_SLICE_X112Y129_AO5),
.O6(CLBLM_L_X74Y129_SLICE_X112Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X74Y129_SLICE_X112Y129_MUXF7A (
.I0(CLBLM_L_X74Y129_SLICE_X112Y129_BO6),
.I1(CLBLM_L_X74Y129_SLICE_X112Y129_AO6),
.O(CLBLM_L_X74Y129_SLICE_X112Y129_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X113Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X113Y129_DO5),
.O6(CLBLM_L_X74Y129_SLICE_X113Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X113Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X113Y129_CO5),
.O6(CLBLM_L_X74Y129_SLICE_X113Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X113Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X113Y129_BO5),
.O6(CLBLM_L_X74Y129_SLICE_X113Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X74Y129_SLICE_X113Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X74Y129_SLICE_X113Y129_AO5),
.O6(CLBLM_L_X74Y129_SLICE_X113Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeae5e04f4a4540)
  ) CLBLM_L_X76Y120_SLICE_X116Y120_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y122_SLICE_X118Y122_DO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_BO6),
.I4(CLBLM_L_X78Y122_SLICE_X120Y122_AO6),
.I5(CLBLL_R_X79Y124_SLICE_X122Y124_CO6),
.O5(CLBLM_L_X76Y120_SLICE_X116Y120_DO5),
.O6(CLBLM_L_X76Y120_SLICE_X116Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbd9eac873516240)
  ) CLBLM_L_X76Y120_SLICE_X116Y120_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLL_R_X77Y114_SLICE_X118Y114_AO6),
.I3(CLBLM_L_X78Y122_SLICE_X120Y122_BO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_DO6),
.I5(CLBLM_L_X78Y123_SLICE_X120Y123_CO6),
.O5(CLBLM_L_X76Y120_SLICE_X116Y120_CO5),
.O6(CLBLM_L_X76Y120_SLICE_X116Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3bbf388c0bbc088)
  ) CLBLM_L_X76Y120_SLICE_X116Y120_BLUT (
.I0(CLBLM_L_X78Y124_SLICE_X120Y124_AO6),
.I1(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I2(CLBLM_L_X78Y123_SLICE_X120Y123_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLM_L_X78Y123_SLICE_X120Y123_AO6),
.I5(CLBLL_R_X77Y129_SLICE_X118Y129_CO6),
.O5(CLBLM_L_X76Y120_SLICE_X116Y120_BO5),
.O6(CLBLM_L_X76Y120_SLICE_X116Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacffac0facf0ac00)
  ) CLBLM_L_X76Y120_SLICE_X116Y120_ALUT (
.I0(CLBLL_R_X77Y122_SLICE_X118Y122_CO6),
.I1(CLBLL_R_X77Y114_SLICE_X118Y114_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y122_SLICE_X118Y122_AO6),
.I5(CLBLM_L_X78Y126_SLICE_X120Y126_BO6),
.O5(CLBLM_L_X76Y120_SLICE_X116Y120_AO5),
.O6(CLBLM_L_X76Y120_SLICE_X116Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y120_SLICE_X116Y120_MUXF7A (
.I0(CLBLM_L_X76Y120_SLICE_X116Y120_BO6),
.I1(CLBLM_L_X76Y120_SLICE_X116Y120_AO6),
.O(CLBLM_L_X76Y120_SLICE_X116Y120_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y120_SLICE_X116Y120_MUXF7B (
.I0(CLBLM_L_X76Y120_SLICE_X116Y120_DO6),
.I1(CLBLM_L_X76Y120_SLICE_X116Y120_CO6),
.O(CLBLM_L_X76Y120_SLICE_X116Y120_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X76Y120_SLICE_X116Y120_MUXF8 (
.I0(CLBLM_L_X76Y120_SLICE_X116Y120_F7BMUX_O),
.I1(CLBLM_L_X76Y120_SLICE_X116Y120_F7AMUX_O),
.O(CLBLM_L_X76Y120_SLICE_X116Y120_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y120_SLICE_X117Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y120_SLICE_X117Y120_DO5),
.O6(CLBLM_L_X76Y120_SLICE_X117Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y120_SLICE_X117Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y120_SLICE_X117Y120_CO5),
.O6(CLBLM_L_X76Y120_SLICE_X117Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y120_SLICE_X117Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y120_SLICE_X117Y120_BO5),
.O6(CLBLM_L_X76Y120_SLICE_X117Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y120_SLICE_X117Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y120_SLICE_X117Y120_AO5),
.O6(CLBLM_L_X76Y120_SLICE_X117Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ffaa5500)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_DLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I4(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_L_X76Y124_SLICE_X116Y124_DO5),
.O6(CLBLM_L_X76Y124_SLICE_X116Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe76dc54ba329810)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I2(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I5(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.O5(CLBLM_L_X76Y124_SLICE_X116Y124_CO5),
.O6(CLBLM_L_X76Y124_SLICE_X116Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222f3c0f3c0)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_BLUT (
.I0(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I4(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X76Y124_SLICE_X116Y124_BO5),
.O6(CLBLM_L_X76Y124_SLICE_X116Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0acac0f00acac)
  ) CLBLM_L_X76Y124_SLICE_X116Y124_ALUT (
.I0(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.O5(CLBLM_L_X76Y124_SLICE_X116Y124_AO5),
.O6(CLBLM_L_X76Y124_SLICE_X116Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y124_SLICE_X116Y124_MUXF7A (
.I0(CLBLM_L_X76Y124_SLICE_X116Y124_BO6),
.I1(CLBLM_L_X76Y124_SLICE_X116Y124_AO6),
.O(CLBLM_L_X76Y124_SLICE_X116Y124_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y124_SLICE_X116Y124_MUXF7B (
.I0(CLBLM_L_X76Y124_SLICE_X116Y124_DO6),
.I1(CLBLM_L_X76Y124_SLICE_X116Y124_CO6),
.O(CLBLM_L_X76Y124_SLICE_X116Y124_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y124_SLICE_X117Y124_DO5),
.O6(CLBLM_L_X76Y124_SLICE_X117Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y124_SLICE_X117Y124_CO5),
.O6(CLBLM_L_X76Y124_SLICE_X117Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y124_SLICE_X117Y124_BO5),
.O6(CLBLM_L_X76Y124_SLICE_X117Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y124_SLICE_X117Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y124_SLICE_X117Y124_AO5),
.O6(CLBLM_L_X76Y124_SLICE_X117Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeae5e04f4a4540)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_DLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I4(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I5(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.O5(CLBLM_L_X76Y125_SLICE_X116Y125_DO5),
.O6(CLBLM_L_X76Y125_SLICE_X116Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4ffe455e4aae400)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_CO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLM_L_X76Y131_SLICE_X116Y131_BO6),
.I5(CLBLM_L_X76Y131_SLICE_X116Y131_AO6),
.O5(CLBLM_L_X76Y125_SLICE_X116Y125_CO5),
.O6(CLBLM_L_X76Y125_SLICE_X116Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf85d58ada80d08)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_BLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_BO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_BO6),
.I4(CLBLL_R_X77Y129_SLICE_X118Y129_AO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_BO6),
.O5(CLBLM_L_X76Y125_SLICE_X116Y125_BO5),
.O6(CLBLM_L_X76Y125_SLICE_X116Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefea4f4ae5e04540)
  ) CLBLM_L_X76Y125_SLICE_X116Y125_ALUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.I4(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I5(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.O5(CLBLM_L_X76Y125_SLICE_X116Y125_AO5),
.O6(CLBLM_L_X76Y125_SLICE_X116Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y125_SLICE_X116Y125_MUXF7A (
.I0(CLBLM_L_X76Y125_SLICE_X116Y125_BO6),
.I1(CLBLM_L_X76Y125_SLICE_X116Y125_AO6),
.O(CLBLM_L_X76Y125_SLICE_X116Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y125_SLICE_X116Y125_MUXF7B (
.I0(CLBLM_L_X76Y125_SLICE_X116Y125_DO6),
.I1(CLBLM_L_X76Y125_SLICE_X116Y125_CO6),
.O(CLBLM_L_X76Y125_SLICE_X116Y125_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X76Y125_SLICE_X116Y125_MUXF8 (
.I0(CLBLM_L_X76Y125_SLICE_X116Y125_F7BMUX_O),
.I1(CLBLM_L_X76Y125_SLICE_X116Y125_F7AMUX_O),
.O(CLBLM_L_X76Y125_SLICE_X116Y125_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacafff0caca0f00)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_DLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I1(CLBLM_L_X98Y132_SLICE_X154Y132_AO6),
.I2(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I3(CLBLM_L_X78Y117_SLICE_X120Y117_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.O5(CLBLM_L_X76Y125_SLICE_X117Y125_DO5),
.O6(CLBLM_L_X76Y125_SLICE_X117Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe455e4aae400e4)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_CLUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I3(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I5(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.O5(CLBLM_L_X76Y125_SLICE_X117Y125_CO5),
.O6(CLBLM_L_X76Y125_SLICE_X117Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0ddddf5a08888)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_BLUT (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.I1(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I2(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I3(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.O5(CLBLM_L_X76Y125_SLICE_X117Y125_BO5),
.O6(CLBLM_L_X76Y125_SLICE_X117Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ff55aa00)
  ) CLBLM_L_X76Y125_SLICE_X117Y125_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I3(CLBLL_R_X79Y125_SLICE_X122Y125_AO6),
.I4(CLBLL_R_X77Y113_SLICE_X118Y113_AO6),
.I5(CLBLM_L_X76Y127_SLICE_X116Y127_CO6),
.O5(CLBLM_L_X76Y125_SLICE_X117Y125_AO5),
.O6(CLBLM_L_X76Y125_SLICE_X117Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y125_SLICE_X117Y125_MUXF7A (
.I0(CLBLM_L_X76Y125_SLICE_X117Y125_BO6),
.I1(CLBLM_L_X76Y125_SLICE_X117Y125_AO6),
.O(CLBLM_L_X76Y125_SLICE_X117Y125_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y125_SLICE_X117Y125_MUXF7B (
.I0(CLBLM_L_X76Y125_SLICE_X117Y125_DO6),
.I1(CLBLM_L_X76Y125_SLICE_X117Y125_CO6),
.O(CLBLM_L_X76Y125_SLICE_X117Y125_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X76Y125_SLICE_X117Y125_MUXF8 (
.I0(CLBLM_L_X76Y125_SLICE_X117Y125_F7BMUX_O),
.I1(CLBLM_L_X76Y125_SLICE_X117Y125_F7AMUX_O),
.O(CLBLM_L_X76Y125_SLICE_X117Y125_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X116Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X116Y127_DO5),
.O6(CLBLM_L_X76Y127_SLICE_X116Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000ff00ff0)
  ) CLBLM_L_X76Y127_SLICE_X116Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(1'b1),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLM_L_X76Y127_SLICE_X116Y127_CO5),
.O6(CLBLM_L_X76Y127_SLICE_X116Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd5df858ad0da808)
  ) CLBLM_L_X76Y127_SLICE_X116Y127_BLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.I4(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.O5(CLBLM_L_X76Y127_SLICE_X116Y127_BO5),
.O6(CLBLM_L_X76Y127_SLICE_X116Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaef4a45e0e5404)
  ) CLBLM_L_X76Y127_SLICE_X116Y127_ALUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.I5(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.O5(CLBLM_L_X76Y127_SLICE_X116Y127_AO5),
.O6(CLBLM_L_X76Y127_SLICE_X116Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y127_SLICE_X116Y127_MUXF7A (
.I0(CLBLM_L_X76Y127_SLICE_X116Y127_BO6),
.I1(CLBLM_L_X76Y127_SLICE_X116Y127_AO6),
.O(CLBLM_L_X76Y127_SLICE_X116Y127_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X117Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X117Y127_DO5),
.O6(CLBLM_L_X76Y127_SLICE_X117Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X117Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X117Y127_CO5),
.O6(CLBLM_L_X76Y127_SLICE_X117Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X117Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X117Y127_BO5),
.O6(CLBLM_L_X76Y127_SLICE_X117Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y127_SLICE_X117Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y127_SLICE_X117Y127_AO5),
.O6(CLBLM_L_X76Y127_SLICE_X117Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3eef322c0eec022)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_DLUT (
.I0(CLBLM_L_X76Y133_SLICE_X117Y133_AO6),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLL_R_X77Y131_SLICE_X118Y131_DO6),
.I3(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I4(CLBLL_R_X77Y131_SLICE_X118Y131_AO6),
.I5(CLBLL_R_X77Y130_SLICE_X118Y130_AO6),
.O5(CLBLM_L_X76Y128_SLICE_X116Y128_DO5),
.O6(CLBLM_L_X76Y128_SLICE_X116Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacaff0fcacaf000)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_CLUT (
.I0(CLBLL_R_X79Y124_SLICE_X122Y124_AO6),
.I1(CLBLM_L_X98Y131_SLICE_X154Y131_AO6),
.I2(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I3(CLBLM_L_X78Y119_SLICE_X120Y119_BO6),
.I4(LIOB33_X0Y79_IOB_X0Y79_I),
.I5(CLBLM_L_X78Y119_SLICE_X120Y119_CO6),
.O5(CLBLM_L_X76Y128_SLICE_X116Y128_CO5),
.O6(CLBLM_L_X76Y128_SLICE_X116Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5eef544a0eea044)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_BLUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLL_R_X77Y133_SLICE_X118Y133_BO6),
.I2(CLBLL_R_X77Y130_SLICE_X118Y130_DO6),
.I3(LIOB33_X0Y79_IOB_X0Y79_I),
.I4(CLBLL_R_X77Y133_SLICE_X118Y133_AO6),
.I5(CLBLL_R_X77Y131_SLICE_X118Y131_CO6),
.O5(CLBLM_L_X76Y128_SLICE_X116Y128_BO5),
.O6(CLBLM_L_X76Y128_SLICE_X116Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfd58f85dad08a80)
  ) CLBLM_L_X76Y128_SLICE_X116Y128_ALUT (
.I0(CLBLL_R_X75Y118_SLICE_X114Y118_DO6),
.I1(CLBLM_L_X78Y129_SLICE_X120Y129_AO6),
.I2(LIOB33_X0Y79_IOB_X0Y79_I),
.I3(CLBLM_L_X78Y120_SLICE_X120Y120_AO6),
.I4(CLBLL_R_X79Y123_SLICE_X122Y123_AO6),
.I5(CLBLM_L_X78Y120_SLICE_X120Y120_BO6),
.O5(CLBLM_L_X76Y128_SLICE_X116Y128_AO5),
.O6(CLBLM_L_X76Y128_SLICE_X116Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7AMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y128_SLICE_X116Y128_MUXF7A (
.I0(CLBLM_L_X76Y128_SLICE_X116Y128_BO6),
.I1(CLBLM_L_X76Y128_SLICE_X116Y128_AO6),
.O(CLBLM_L_X76Y128_SLICE_X116Y128_F7AMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F7BMUX" *)
  MUXF7 #(
  ) CLBLM_L_X76Y128_SLICE_X116Y128_MUXF7B (
.I0(CLBLM_L_X76Y128_SLICE_X116Y128_DO6),
.I1(CLBLM_L_X76Y128_SLICE_X116Y128_CO6),
.O(CLBLM_L_X76Y128_SLICE_X116Y128_F7BMUX_O),
.S(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "F8MUX" *)
  MUXF8 #(
  ) CLBLM_L_X76Y128_SLICE_X116Y128_MUXF8 (
.I0(CLBLM_L_X76Y128_SLICE_X116Y128_F7BMUX_O),
.I1(CLBLM_L_X76Y128_SLICE_X116Y128_F7AMUX_O),
.O(CLBLM_L_X76Y128_SLICE_X116Y128_F8MUX_O),
.S(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y128_SLICE_X117Y128_DO5),
.O6(CLBLM_L_X76Y128_SLICE_X117Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y128_SLICE_X117Y128_CO5),
.O6(CLBLM_L_X76Y128_SLICE_X117Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y128_SLICE_X117Y128_BO5),
.O6(CLBLM_L_X76Y128_SLICE_X117Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y128_SLICE_X117Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y128_SLICE_X117Y128_AO5),
.O6(CLBLM_L_X76Y128_SLICE_X117Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y131_SLICE_X116Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y131_SLICE_X116Y131_DO5),
.O6(CLBLM_L_X76Y131_SLICE_X116Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y131_SLICE_X116Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y131_SLICE_X116Y131_CO5),
.O6(CLBLM_L_X76Y131_SLICE_X116Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeae5404efea4540)
  ) CLBLM_L_X76Y131_SLICE_X116Y131_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(RIOB33_X105Y147_IOB_X1Y148_I),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(LIOB33_X0Y197_IOB_X0Y198_I),
.I4(RIOB33_X105Y91_IOB_X1Y92_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLM_L_X76Y131_SLICE_X116Y131_BO5),
.O6(CLBLM_L_X76Y131_SLICE_X116Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb51ea40fe54ba10)
  ) CLBLM_L_X76Y131_SLICE_X116Y131_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(LIOB33_X0Y183_IOB_X0Y184_I),
.I3(RIOB33_X105Y77_IOB_X1Y78_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLM_L_X76Y131_SLICE_X116Y131_AO5),
.O6(CLBLM_L_X76Y131_SLICE_X116Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y131_SLICE_X117Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y131_SLICE_X117Y131_DO5),
.O6(CLBLM_L_X76Y131_SLICE_X117Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y131_SLICE_X117Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y131_SLICE_X117Y131_CO5),
.O6(CLBLM_L_X76Y131_SLICE_X117Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y131_SLICE_X117Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y131_SLICE_X117Y131_BO5),
.O6(CLBLM_L_X76Y131_SLICE_X117Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y131_SLICE_X117Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y131_SLICE_X117Y131_AO5),
.O6(CLBLM_L_X76Y131_SLICE_X117Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X116Y133_DO5),
.O6(CLBLM_L_X76Y133_SLICE_X116Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X116Y133_CO5),
.O6(CLBLM_L_X76Y133_SLICE_X116Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X116Y133_BO5),
.O6(CLBLM_L_X76Y133_SLICE_X116Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X116Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X116Y133_AO5),
.O6(CLBLM_L_X76Y133_SLICE_X116Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X117Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X117Y133_DO5),
.O6(CLBLM_L_X76Y133_SLICE_X117Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X117Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X117Y133_CO5),
.O6(CLBLM_L_X76Y133_SLICE_X117Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X76Y133_SLICE_X117Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X76Y133_SLICE_X117Y133_BO5),
.O6(CLBLM_L_X76Y133_SLICE_X117Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5a0f5a0e4e4)
  ) CLBLM_L_X76Y133_SLICE_X117Y133_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(LIOB33_X0Y189_IOB_X0Y190_I),
.I2(RIOB33_X105Y83_IOB_X1Y84_I),
.I3(RIOB33_X105Y139_IOB_X1Y140_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLM_L_X76Y133_SLICE_X117Y133_AO5),
.O6(CLBLM_L_X76Y133_SLICE_X117Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y117_SLICE_X120Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y117_SLICE_X120Y117_DO5),
.O6(CLBLM_L_X78Y117_SLICE_X120Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y117_SLICE_X120Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y117_SLICE_X120Y117_CO5),
.O6(CLBLM_L_X78Y117_SLICE_X120Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc5acca5cc00)
  ) CLBLM_L_X78Y117_SLICE_X120Y117_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(LIOB33_X0Y155_IOB_X0Y155_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_L_X78Y117_SLICE_X120Y117_BO5),
.O6(CLBLM_L_X78Y117_SLICE_X120Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4d8d8)
  ) CLBLM_L_X78Y117_SLICE_X120Y117_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y117_IOB_X1Y117_I),
.I2(LIOB33_X0Y161_IOB_X0Y161_I),
.I3(RIOB33_X105Y55_IOB_X1Y55_I),
.I4(LIOB33_X0Y85_IOB_X0Y85_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLM_L_X78Y117_SLICE_X120Y117_AO5),
.O6(CLBLM_L_X78Y117_SLICE_X120Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y117_SLICE_X121Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y117_SLICE_X121Y117_DO5),
.O6(CLBLM_L_X78Y117_SLICE_X121Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y117_SLICE_X121Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y117_SLICE_X121Y117_CO5),
.O6(CLBLM_L_X78Y117_SLICE_X121Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y117_SLICE_X121Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y117_SLICE_X121Y117_BO5),
.O6(CLBLM_L_X78Y117_SLICE_X121Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y117_SLICE_X121Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y117_SLICE_X121Y117_AO5),
.O6(CLBLM_L_X78Y117_SLICE_X121Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y119_SLICE_X120Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y119_SLICE_X120Y119_DO5),
.O6(CLBLM_L_X78Y119_SLICE_X120Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffc33c00)
  ) CLBLM_L_X78Y119_SLICE_X120Y119_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(LIOB33_X0Y83_IOB_X0Y84_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y153_IOB_X0Y154_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLM_L_X78Y119_SLICE_X120Y119_CO5),
.O6(CLBLM_L_X78Y119_SLICE_X120Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffed00edff480048)
  ) CLBLM_L_X78Y119_SLICE_X120Y119_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(RIOB33_X105Y55_IOB_X1Y56_I),
.I5(LIOB33_X0Y161_IOB_X0Y162_I),
.O5(CLBLM_L_X78Y119_SLICE_X120Y119_BO5),
.O6(CLBLM_L_X78Y119_SLICE_X120Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdec3120fedc3210)
  ) CLBLM_L_X78Y119_SLICE_X120Y119_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(LIOB33_X0Y159_IOB_X0Y160_I),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(RIOB33_X105Y53_IOB_X1Y54_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLM_L_X78Y119_SLICE_X120Y119_AO5),
.O6(CLBLM_L_X78Y119_SLICE_X120Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y119_SLICE_X121Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y119_SLICE_X121Y119_DO5),
.O6(CLBLM_L_X78Y119_SLICE_X121Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y119_SLICE_X121Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y119_SLICE_X121Y119_CO5),
.O6(CLBLM_L_X78Y119_SLICE_X121Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y119_SLICE_X121Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y119_SLICE_X121Y119_BO5),
.O6(CLBLM_L_X78Y119_SLICE_X121Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y119_SLICE_X121Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y119_SLICE_X121Y119_AO5),
.O6(CLBLM_L_X78Y119_SLICE_X121Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X120Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X120Y120_DO5),
.O6(CLBLM_L_X78Y120_SLICE_X120Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000be82be82)
  ) CLBLM_L_X78Y120_SLICE_X120Y120_CLUT (
.I0(LIOB33_X0Y163_IOB_X0Y164_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(RIOB33_X105Y119_IOB_X1Y120_I),
.I4(RIOB33_X105Y57_IOB_X1Y58_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLM_L_X78Y120_SLICE_X120Y120_CO5),
.O6(CLBLM_L_X78Y120_SLICE_X120Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5cca0ccfacc50)
  ) CLBLM_L_X78Y120_SLICE_X120Y120_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y153_IOB_X0Y153_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLM_L_X78Y120_SLICE_X120Y120_BO5),
.O6(CLBLM_L_X78Y120_SLICE_X120Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff900f9ff600060)
  ) CLBLM_L_X78Y120_SLICE_X120Y120_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(LIOB33_X0Y83_IOB_X0Y83_I),
.I4(RIOB33_X105Y57_IOB_X1Y57_I),
.I5(LIOB33_X0Y163_IOB_X0Y163_I),
.O5(CLBLM_L_X78Y120_SLICE_X120Y120_AO5),
.O6(CLBLM_L_X78Y120_SLICE_X120Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X121Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X121Y120_DO5),
.O6(CLBLM_L_X78Y120_SLICE_X121Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X121Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X121Y120_CO5),
.O6(CLBLM_L_X78Y120_SLICE_X121Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X121Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X121Y120_BO5),
.O6(CLBLM_L_X78Y120_SLICE_X121Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y120_SLICE_X121Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y120_SLICE_X121Y120_AO5),
.O6(CLBLM_L_X78Y120_SLICE_X121Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X120Y121_DO5),
.O6(CLBLM_L_X78Y121_SLICE_X120Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X120Y121_CO5),
.O6(CLBLM_L_X78Y121_SLICE_X120Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X120Y121_BO5),
.O6(CLBLM_L_X78Y121_SLICE_X120Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31fe32ec20dc10)
  ) CLBLM_L_X78Y121_SLICE_X120Y121_ALUT (
.I0(LIOB33_X0Y85_IOB_X0Y85_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(LIOB33_X0Y165_IOB_X0Y165_I),
.I3(RIOB33_X105Y59_IOB_X1Y59_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X78Y121_SLICE_X120Y121_AO5),
.O6(CLBLM_L_X78Y121_SLICE_X120Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X121Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X121Y121_DO5),
.O6(CLBLM_L_X78Y121_SLICE_X121Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X121Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X121Y121_CO5),
.O6(CLBLM_L_X78Y121_SLICE_X121Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X121Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X121Y121_BO5),
.O6(CLBLM_L_X78Y121_SLICE_X121Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y121_SLICE_X121Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y121_SLICE_X121Y121_AO5),
.O6(CLBLM_L_X78Y121_SLICE_X121Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y122_SLICE_X120Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y122_SLICE_X120Y122_DO5),
.O6(CLBLM_L_X78Y122_SLICE_X120Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y122_SLICE_X120Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y122_SLICE_X120Y122_CO5),
.O6(CLBLM_L_X78Y122_SLICE_X120Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5facccca050)
  ) CLBLM_L_X78Y122_SLICE_X120Y122_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y59_IOB_X1Y60_I),
.I2(LIOB33_X0Y165_IOB_X0Y166_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(LIOB33_X0Y83_IOB_X0Y83_I),
.I5(RIOB33_X105Y121_IOB_X1Y122_I),
.O5(CLBLM_L_X78Y122_SLICE_X120Y122_BO5),
.O6(CLBLM_L_X78Y122_SLICE_X120Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ee44f0f0dd88)
  ) CLBLM_L_X78Y122_SLICE_X120Y122_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(RIOB33_X105Y87_IOB_X1Y87_I),
.I3(LIOB33_X0Y193_IOB_X0Y193_I),
.I4(LIOB33_X0Y83_IOB_X0Y83_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLM_L_X78Y122_SLICE_X120Y122_AO5),
.O6(CLBLM_L_X78Y122_SLICE_X120Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y122_SLICE_X121Y122_DO5),
.O6(CLBLM_L_X78Y122_SLICE_X121Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y122_SLICE_X121Y122_CO5),
.O6(CLBLM_L_X78Y122_SLICE_X121Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y122_SLICE_X121Y122_BO5),
.O6(CLBLM_L_X78Y122_SLICE_X121Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y122_SLICE_X121Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y122_SLICE_X121Y122_AO5),
.O6(CLBLM_L_X78Y122_SLICE_X121Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000accaacca)
  ) CLBLM_L_X78Y123_SLICE_X120Y123_DLUT (
.I0(LIOB33_X0Y171_IOB_X0Y171_I),
.I1(RIOB33_X105Y125_IOB_X1Y126_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(RIOB33_X105Y65_IOB_X1Y65_I),
.I5(LIOB33_X0Y83_IOB_X0Y83_I),
.O5(CLBLM_L_X78Y123_SLICE_X120Y123_DO5),
.O6(CLBLM_L_X78Y123_SLICE_X120Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeafeae45405404)
  ) CLBLM_L_X78Y123_SLICE_X120Y123_CLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(LIOB33_SING_X0Y199_IOB_X0Y199_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(RIOB33_X105Y93_IOB_X1Y93_I),
.O5(CLBLM_L_X78Y123_SLICE_X120Y123_CO5),
.O6(CLBLM_L_X78Y123_SLICE_X120Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefd0e0df4f80408)
  ) CLBLM_L_X78Y123_SLICE_X120Y123_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(RIOB33_X105Y85_IOB_X1Y86_I),
.I5(LIOB33_X0Y191_IOB_X0Y192_I),
.O5(CLBLM_L_X78Y123_SLICE_X120Y123_BO5),
.O6(CLBLM_L_X78Y123_SLICE_X120Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefd0e0df4f80408)
  ) CLBLM_L_X78Y123_SLICE_X120Y123_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y189_IOB_X1Y190_I),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(RIOB33_X105Y73_IOB_X1Y74_I),
.I5(LIOB33_X0Y179_IOB_X0Y180_I),
.O5(CLBLM_L_X78Y123_SLICE_X120Y123_AO5),
.O6(CLBLM_L_X78Y123_SLICE_X120Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y123_SLICE_X121Y123_DO5),
.O6(CLBLM_L_X78Y123_SLICE_X121Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y123_SLICE_X121Y123_CO5),
.O6(CLBLM_L_X78Y123_SLICE_X121Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y123_SLICE_X121Y123_BO5),
.O6(CLBLM_L_X78Y123_SLICE_X121Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y123_SLICE_X121Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y123_SLICE_X121Y123_AO5),
.O6(CLBLM_L_X78Y123_SLICE_X121Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X120Y124_DO5),
.O6(CLBLM_L_X78Y124_SLICE_X120Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X120Y124_CO5),
.O6(CLBLM_L_X78Y124_SLICE_X120Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc5cacac5c0c0)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(RIOB33_X105Y81_IOB_X1Y82_I),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(LIOB33_X0Y85_IOB_X0Y85_I),
.I4(LIOB33_X0Y187_IOB_X0Y188_I),
.I5(RIOB33_X105Y137_IOB_X1Y138_I),
.O5(CLBLM_L_X78Y124_SLICE_X120Y124_BO5),
.O6(CLBLM_L_X78Y124_SLICE_X120Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfedc3210fdec3120)
  ) CLBLM_L_X78Y124_SLICE_X120Y124_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y84_I),
.I1(LIOB33_X0Y83_IOB_X0Y83_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(LIOB33_X0Y185_IOB_X0Y185_I),
.I4(RIOB33_X105Y79_IOB_X1Y79_I),
.I5(LIOB33_X0Y85_IOB_X0Y85_I),
.O5(CLBLM_L_X78Y124_SLICE_X120Y124_AO5),
.O6(CLBLM_L_X78Y124_SLICE_X120Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X121Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X121Y124_DO5),
.O6(CLBLM_L_X78Y124_SLICE_X121Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X121Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X121Y124_CO5),
.O6(CLBLM_L_X78Y124_SLICE_X121Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X121Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X121Y124_BO5),
.O6(CLBLM_L_X78Y124_SLICE_X121Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y124_SLICE_X121Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y124_SLICE_X121Y124_AO5),
.O6(CLBLM_L_X78Y124_SLICE_X121Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y126_SLICE_X120Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y126_SLICE_X120Y126_DO5),
.O6(CLBLM_L_X78Y126_SLICE_X120Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y126_SLICE_X120Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y126_SLICE_X120Y126_CO5),
.O6(CLBLM_L_X78Y126_SLICE_X120Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0df808fe0ef404)
  ) CLBLM_L_X78Y126_SLICE_X120Y126_BLUT (
.I0(LIOB33_X0Y85_IOB_X0Y85_I),
.I1(LIOB33_X0Y181_IOB_X0Y181_I),
.I2(LIOB33_X0Y83_IOB_X0Y83_I),
.I3(RIOB33_X105Y75_IOB_X1Y75_I),
.I4(RIOB33_X105Y191_IOB_X1Y191_I),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLM_L_X78Y126_SLICE_X120Y126_BO5),
.O6(CLBLM_L_X78Y126_SLICE_X120Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e4e4ff00d8d8)
  ) CLBLM_L_X78Y126_SLICE_X120Y126_ALUT (
.I0(LIOB33_X0Y85_IOB_X0Y85_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(LIOB33_X0Y187_IOB_X0Y187_I),
.I3(RIOB33_X105Y81_IOB_X1Y81_I),
.I4(LIOB33_X0Y83_IOB_X0Y83_I),
.I5(LIOB33_X0Y83_IOB_X0Y84_I),
.O5(CLBLM_L_X78Y126_SLICE_X120Y126_AO5),
.O6(CLBLM_L_X78Y126_SLICE_X120Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y126_SLICE_X121Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y126_SLICE_X121Y126_DO5),
.O6(CLBLM_L_X78Y126_SLICE_X121Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y126_SLICE_X121Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y126_SLICE_X121Y126_CO5),
.O6(CLBLM_L_X78Y126_SLICE_X121Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y126_SLICE_X121Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y126_SLICE_X121Y126_BO5),
.O6(CLBLM_L_X78Y126_SLICE_X121Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y126_SLICE_X121Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y126_SLICE_X121Y126_AO5),
.O6(CLBLM_L_X78Y126_SLICE_X121Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X120Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X120Y129_DO5),
.O6(CLBLM_L_X78Y129_SLICE_X120Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X120Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X120Y129_CO5),
.O6(CLBLM_L_X78Y129_SLICE_X120Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X120Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X120Y129_BO5),
.O6(CLBLM_L_X78Y129_SLICE_X120Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfe5154eaba4010)
  ) CLBLM_L_X78Y129_SLICE_X120Y129_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(LIOB33_X0Y85_IOB_X0Y85_I),
.I2(LIOB33_X0Y173_IOB_X0Y174_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(RIOB33_X105Y67_IOB_X1Y68_I),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_L_X78Y129_SLICE_X120Y129_AO5),
.O6(CLBLM_L_X78Y129_SLICE_X120Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X121Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X121Y129_DO5),
.O6(CLBLM_L_X78Y129_SLICE_X121Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X121Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X121Y129_CO5),
.O6(CLBLM_L_X78Y129_SLICE_X121Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X121Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X121Y129_BO5),
.O6(CLBLM_L_X78Y129_SLICE_X121Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X78Y129_SLICE_X121Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X78Y129_SLICE_X121Y129_AO5),
.O6(CLBLM_L_X78Y129_SLICE_X121Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X154Y131_DO5),
.O6(CLBLM_L_X98Y131_SLICE_X154Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X154Y131_CO5),
.O6(CLBLM_L_X98Y131_SLICE_X154Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X154Y131_BO5),
.O6(CLBLM_L_X98Y131_SLICE_X154Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefafaee44505044)
  ) CLBLM_L_X98Y131_SLICE_X154Y131_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(RIOB33_X105Y187_IOB_X1Y187_I),
.I2(RIOB33_SING_X105Y199_IOB_X1Y199_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(LIOB33_X0Y85_IOB_X0Y85_I),
.I5(RIOB33_SING_X105Y99_IOB_X1Y99_I),
.O5(CLBLM_L_X98Y131_SLICE_X154Y131_AO5),
.O6(CLBLM_L_X98Y131_SLICE_X154Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X155Y131_DO5),
.O6(CLBLM_L_X98Y131_SLICE_X155Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X155Y131_CO5),
.O6(CLBLM_L_X98Y131_SLICE_X155Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X155Y131_BO5),
.O6(CLBLM_L_X98Y131_SLICE_X155Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y131_SLICE_X155Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y131_SLICE_X155Y131_AO5),
.O6(CLBLM_L_X98Y131_SLICE_X155Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X154Y132_DO5),
.O6(CLBLM_L_X98Y132_SLICE_X154Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X154Y132_CO5),
.O6(CLBLM_L_X98Y132_SLICE_X154Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X154Y132_BO5),
.O6(CLBLM_L_X98Y132_SLICE_X154Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffebbeaa55411400)
  ) CLBLM_L_X98Y132_SLICE_X154Y132_ALUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(LIOB33_X0Y83_IOB_X0Y84_I),
.I2(LIOB33_X0Y85_IOB_X0Y85_I),
.I3(RIOB33_X105Y197_IOB_X1Y198_I),
.I4(RIOB33_X105Y185_IOB_X1Y186_I),
.I5(RIOB33_X105Y97_IOB_X1Y98_I),
.O5(CLBLM_L_X98Y132_SLICE_X154Y132_AO5),
.O6(CLBLM_L_X98Y132_SLICE_X154Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X155Y132_DO5),
.O6(CLBLM_L_X98Y132_SLICE_X155Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X155Y132_CO5),
.O6(CLBLM_L_X98Y132_SLICE_X155Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X155Y132_BO5),
.O6(CLBLM_L_X98Y132_SLICE_X155Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X98Y132_SLICE_X155Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X98Y132_SLICE_X155Y132_AO5),
.O6(CLBLM_L_X98Y132_SLICE_X155Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y120_SLICE_X0Y120_DO6),
.Q(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001fefffffe0100)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_CO6),
.I4(CLBLL_L_X2Y123_SLICE_X0Y123_BQ),
.I5(CLBLL_R_X71Y125_SLICE_X106Y125_DO6),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333336ccccc9cc)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(CLBLL_R_X71Y125_SLICE_X106Y125_CO6),
.I2(LIOB33_X0Y81_IOB_X0Y81_I),
.I3(CLBLL_L_X2Y123_SLICE_X1Y123_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y82_I),
.I5(CLBLL_L_X2Y124_SLICE_X0Y124_AQ),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y116_SLICE_X74Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y116_SLICE_X74Y116_DO5),
.O6(CLBLM_R_X49Y116_SLICE_X74Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y116_SLICE_X74Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y116_SLICE_X74Y116_CO5),
.O6(CLBLM_R_X49Y116_SLICE_X74Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y116_SLICE_X74Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y116_SLICE_X74Y116_BO5),
.O6(CLBLM_R_X49Y116_SLICE_X74Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X49Y116_SLICE_X74Y116_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(LIOB33_X0Y81_IOB_X0Y81_I),
.I2(LIOB33_X0Y81_IOB_X0Y82_I),
.I3(LIOB33_X0Y83_IOB_X0Y84_I),
.I4(LIOB33_X0Y83_IOB_X0Y83_I),
.I5(LIOB33_X0Y79_IOB_X0Y80_I),
.O5(CLBLM_R_X49Y116_SLICE_X74Y116_AO5),
.O6(CLBLM_R_X49Y116_SLICE_X74Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y116_SLICE_X75Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y116_SLICE_X75Y116_DO5),
.O6(CLBLM_R_X49Y116_SLICE_X75Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y116_SLICE_X75Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y116_SLICE_X75Y116_CO5),
.O6(CLBLM_R_X49Y116_SLICE_X75Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y116_SLICE_X75Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y116_SLICE_X75Y116_BO5),
.O6(CLBLM_R_X49Y116_SLICE_X75Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X49Y116_SLICE_X75Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X49Y116_SLICE_X75Y116_AO5),
.O6(CLBLM_R_X49Y116_SLICE_X75Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y117_SLICE_X88Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_R_X59Y118_SLICE_X88Y118_AO6),
.Q(CLBLM_R_X59Y117_SLICE_X88Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y117_SLICE_X88Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y117_SLICE_X88Y117_DO5),
.O6(CLBLM_R_X59Y117_SLICE_X88Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y117_SLICE_X88Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y117_SLICE_X88Y117_CO5),
.O6(CLBLM_R_X59Y117_SLICE_X88Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y117_SLICE_X88Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y117_SLICE_X88Y117_BO5),
.O6(CLBLM_R_X59Y117_SLICE_X88Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88bb88b8b8)
  ) CLBLM_R_X59Y117_SLICE_X88Y117_ALUT (
.I0(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I1(CLBLM_R_X49Y116_SLICE_X74Y116_AO6),
.I2(CLBLM_R_X59Y117_SLICE_X88Y117_AQ),
.I3(CLBLM_R_X59Y118_SLICE_X88Y118_AQ),
.I4(CLBLM_L_X46Y116_SLICE_X70Y116_AO6),
.I5(CLBLM_L_X46Y116_SLICE_X70Y116_BO6),
.O5(CLBLM_R_X59Y117_SLICE_X88Y117_AO5),
.O6(CLBLM_R_X59Y117_SLICE_X88Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y117_SLICE_X89Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y117_SLICE_X89Y117_DO5),
.O6(CLBLM_R_X59Y117_SLICE_X89Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y117_SLICE_X89Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y117_SLICE_X89Y117_CO5),
.O6(CLBLM_R_X59Y117_SLICE_X89Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y117_SLICE_X89Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y117_SLICE_X89Y117_BO5),
.O6(CLBLM_R_X59Y117_SLICE_X89Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y117_SLICE_X89Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y117_SLICE_X89Y117_AO5),
.O6(CLBLM_R_X59Y117_SLICE_X89Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X59Y118_SLICE_X88Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O),
.CE(1'b1),
.D(CLBLM_R_X59Y117_SLICE_X88Y117_AO6),
.Q(CLBLM_R_X59Y118_SLICE_X88Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y118_SLICE_X88Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y118_SLICE_X88Y118_DO5),
.O6(CLBLM_R_X59Y118_SLICE_X88Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y118_SLICE_X88Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y118_SLICE_X88Y118_CO5),
.O6(CLBLM_R_X59Y118_SLICE_X88Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f5a0ee44)
  ) CLBLM_R_X59Y118_SLICE_X88Y118_BLUT (
.I0(LIOB33_X0Y83_IOB_X0Y83_I),
.I1(RIOB33_X105Y163_IOB_X1Y164_I),
.I2(CLBLM_R_X59Y118_SLICE_X88Y118_AQ),
.I3(CLBLM_R_X59Y117_SLICE_X88Y117_AQ),
.I4(LIOB33_X0Y83_IOB_X0Y84_I),
.I5(CLBLM_L_X44Y118_SLICE_X66Y118_AO6),
.O5(CLBLM_R_X59Y118_SLICE_X88Y118_BO5),
.O6(CLBLM_R_X59Y118_SLICE_X88Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e1ff0f0f1e0)
  ) CLBLM_R_X59Y118_SLICE_X88Y118_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y80_I),
.I1(LIOB33_X0Y81_IOB_X0Y82_I),
.I2(CLBLM_R_X59Y118_SLICE_X88Y118_AQ),
.I3(CLBLM_R_X59Y118_SLICE_X88Y118_BO6),
.I4(LIOB33_X0Y81_IOB_X0Y81_I),
.I5(CLBLL_R_X73Y122_SLICE_X110Y122_BO6),
.O5(CLBLM_R_X59Y118_SLICE_X88Y118_AO5),
.O6(CLBLM_R_X59Y118_SLICE_X88Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y118_SLICE_X89Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y118_SLICE_X89Y118_DO5),
.O6(CLBLM_R_X59Y118_SLICE_X89Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y118_SLICE_X89Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y118_SLICE_X89Y118_CO5),
.O6(CLBLM_R_X59Y118_SLICE_X89Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y118_SLICE_X89Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y118_SLICE_X89Y118_BO5),
.O6(CLBLM_R_X59Y118_SLICE_X89Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X59Y118_SLICE_X89Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X59Y118_SLICE_X89Y118_AO5),
.O6(CLBLM_R_X59Y118_SLICE_X89Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y80_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y80_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y81_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y81_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y81_IOB_X0Y82_IBUF (
.I(LIOB33_X0Y81_IOB_X0Y82_IPAD),
.O(LIOB33_X0Y81_IOB_X0Y82_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y83_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y83_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y83_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y83_IOB_X0Y84_IBUF (
.I(LIOB33_X0Y83_IOB_X0Y84_IPAD),
.O(LIOB33_X0Y83_IOB_X0Y84_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y85_IOB_X0Y85_IBUF (
.I(LIOB33_X0Y85_IOB_X0Y85_IPAD),
.O(LIOB33_X0Y85_IOB_X0Y85_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y85_IOB_X0Y86_OBUF (
.I(CLBLM_L_X70Y119_SLICE_X104Y119_AO6),
.O(LIOB33_X0Y85_IOB_X0Y86_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y87_IOB_X0Y87_OBUF (
.I(CLBLL_R_X71Y119_SLICE_X106Y119_AO6),
.O(LIOB33_X0Y87_IOB_X0Y87_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y87_IOB_X0Y88_OBUF (
.I(CLBLM_L_X70Y128_SLICE_X105Y128_AO6),
.O(LIOB33_X0Y87_IOB_X0Y88_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y89_IOB_X0Y89_OBUF (
.I(CLBLM_L_X70Y128_SLICE_X105Y128_CO6),
.O(LIOB33_X0Y89_IOB_X0Y89_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y89_IOB_X0Y90_OBUF (
.I(CLBLL_R_X71Y128_SLICE_X106Y128_AO6),
.O(LIOB33_X0Y89_IOB_X0Y90_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y91_IOB_X0Y91_OBUF (
.I(CLBLL_R_X71Y128_SLICE_X106Y128_CO6),
.O(LIOB33_X0Y91_IOB_X0Y91_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y91_IOB_X0Y92_OBUF (
.I(CLBLL_R_X71Y131_SLICE_X107Y131_BO6),
.O(LIOB33_X0Y91_IOB_X0Y92_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y93_IOB_X0Y93_OBUF (
.I(CLBLL_R_X71Y131_SLICE_X107Y131_DO6),
.O(LIOB33_X0Y93_IOB_X0Y93_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y93_IOB_X0Y94_OBUF (
.I(CLBLM_L_X70Y129_SLICE_X104Y129_AO6),
.O(LIOB33_X0Y93_IOB_X0Y94_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y95_IOB_X0Y95_OBUF (
.I(CLBLM_L_X70Y129_SLICE_X104Y129_CO6),
.O(LIOB33_X0Y95_IOB_X0Y95_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y95_IOB_X0Y96_OBUF (
.I(CLBLM_L_X70Y124_SLICE_X104Y124_AO6),
.O(LIOB33_X0Y95_IOB_X0Y96_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y97_IOB_X0Y97_OBUF (
.I(CLBLM_L_X70Y124_SLICE_X104Y124_CO6),
.O(LIOB33_X0Y97_IOB_X0Y97_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y97_IOB_X0Y98_OBUF (
.I(CLBLL_R_X71Y131_SLICE_X106Y131_AO6),
.O(LIOB33_X0Y97_IOB_X0Y98_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLM_R_X59Y117_SLICE_X88Y117_AO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y105_SLICE_X0Y105_CO6),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLM_L_X56Y116_SLICE_X84Y116_AO6),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLM_L_X56Y116_SLICE_X84Y116_CO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLM_L_X70Y121_SLICE_X104Y121_AO6),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLM_L_X70Y123_SLICE_X104Y123_BO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_L_X70Y123_SLICE_X105Y123_AO6),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLM_L_X70Y123_SLICE_X105Y123_CO6),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_L_X72Y131_SLICE_X108Y131_AO6),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLL_R_X71Y131_SLICE_X107Y131_AO6),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_L_X70Y122_SLICE_X104Y122_AO6),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_L_X70Y122_SLICE_X104Y122_CO6),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X70Y121_SLICE_X105Y121_AO6),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_L_X70Y121_SLICE_X105Y121_CO6),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_L_X70Y119_SLICE_X105Y119_AO6),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X70Y119_SLICE_X105Y119_CO6),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_L_X70Y121_SLICE_X104Y121_BO6),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X70Y121_SLICE_X104Y121_DO6),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_L_X70Y127_SLICE_X104Y127_AO6),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_L_X70Y128_SLICE_X104Y128_BO6),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_L_X70Y123_SLICE_X105Y123_DO6),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X70Y124_SLICE_X105Y124_BO6),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_L_X70Y127_SLICE_X104Y127_BO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_L_X70Y127_SLICE_X104Y127_DO6),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_CO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLL_L_X2Y124_SLICE_X1Y124_AO6),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X2Y123_SLICE_X1Y123_AO6),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLL_L_X2Y124_SLICE_X0Y124_AO6),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X2Y124_SLICE_X0Y124_CO6),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X2Y124_SLICE_X1Y124_CO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X2Y124_SLICE_X0Y124_DO6),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X2Y123_SLICE_X0Y123_AO6),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X2Y123_SLICE_X0Y123_CO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_DO6),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X2Y119_SLICE_X1Y119_CO6),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X2Y121_SLICE_X0Y121_DO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_L_X2Y123_SLICE_X0Y123_DO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y151_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y151_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y151_IOB_X0Y152_IBUF (
.I(LIOB33_X0Y151_IOB_X0Y152_IPAD),
.O(LIOB33_X0Y151_IOB_X0Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y153_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y153_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y153_IOB_X0Y154_IBUF (
.I(LIOB33_X0Y153_IOB_X0Y154_IPAD),
.O(LIOB33_X0Y153_IOB_X0Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y155_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y155_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y155_IOB_X0Y156_IBUF (
.I(LIOB33_X0Y155_IOB_X0Y156_IPAD),
.O(LIOB33_X0Y155_IOB_X0Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y157_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y157_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y157_IOB_X0Y158_IBUF (
.I(LIOB33_X0Y157_IOB_X0Y158_IPAD),
.O(LIOB33_X0Y157_IOB_X0Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y159_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y159_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y159_IOB_X0Y160_IBUF (
.I(LIOB33_X0Y159_IOB_X0Y160_IPAD),
.O(LIOB33_X0Y159_IOB_X0Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y161_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y161_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y161_IOB_X0Y162_IBUF (
.I(LIOB33_X0Y161_IOB_X0Y162_IPAD),
.O(LIOB33_X0Y161_IOB_X0Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y163_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y163_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y163_IOB_X0Y164_IBUF (
.I(LIOB33_X0Y163_IOB_X0Y164_IPAD),
.O(LIOB33_X0Y163_IOB_X0Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y165_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y165_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y165_IOB_X0Y166_IBUF (
.I(LIOB33_X0Y165_IOB_X0Y166_IPAD),
.O(LIOB33_X0Y165_IOB_X0Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y167_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y167_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y167_IOB_X0Y168_IBUF (
.I(LIOB33_X0Y167_IOB_X0Y168_IPAD),
.O(LIOB33_X0Y167_IOB_X0Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y169_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y169_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y169_IOB_X0Y170_IBUF (
.I(LIOB33_X0Y169_IOB_X0Y170_IPAD),
.O(LIOB33_X0Y169_IOB_X0Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y171_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y171_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y171_IOB_X0Y172_IBUF (
.I(LIOB33_X0Y171_IOB_X0Y172_IPAD),
.O(LIOB33_X0Y171_IOB_X0Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y173_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y173_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y173_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y173_IOB_X0Y174_IBUF (
.I(LIOB33_X0Y173_IOB_X0Y174_IPAD),
.O(LIOB33_X0Y173_IOB_X0Y174_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y175_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y175_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y175_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y175_IOB_X0Y176_IBUF (
.I(LIOB33_X0Y175_IOB_X0Y176_IPAD),
.O(LIOB33_X0Y175_IOB_X0Y176_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y177_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y177_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y177_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y177_IOB_X0Y178_IBUF (
.I(LIOB33_X0Y177_IOB_X0Y178_IPAD),
.O(LIOB33_X0Y177_IOB_X0Y178_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y179_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y179_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y179_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y179_IOB_X0Y180_IBUF (
.I(LIOB33_X0Y179_IOB_X0Y180_IPAD),
.O(LIOB33_X0Y179_IOB_X0Y180_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y181_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y181_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y181_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y181_IOB_X0Y182_IBUF (
.I(LIOB33_X0Y181_IOB_X0Y182_IPAD),
.O(LIOB33_X0Y181_IOB_X0Y182_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y183_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y183_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y183_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y183_IOB_X0Y184_IBUF (
.I(LIOB33_X0Y183_IOB_X0Y184_IPAD),
.O(LIOB33_X0Y183_IOB_X0Y184_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y185_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y185_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y185_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y185_IOB_X0Y186_IBUF (
.I(LIOB33_X0Y185_IOB_X0Y186_IPAD),
.O(LIOB33_X0Y185_IOB_X0Y186_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y187_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y187_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y187_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y187_IOB_X0Y188_IBUF (
.I(LIOB33_X0Y187_IOB_X0Y188_IPAD),
.O(LIOB33_X0Y187_IOB_X0Y188_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y189_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y189_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y189_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y189_IOB_X0Y190_IBUF (
.I(LIOB33_X0Y189_IOB_X0Y190_IPAD),
.O(LIOB33_X0Y189_IOB_X0Y190_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y191_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y191_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y191_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y191_IOB_X0Y192_IBUF (
.I(LIOB33_X0Y191_IOB_X0Y192_IPAD),
.O(LIOB33_X0Y191_IOB_X0Y192_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y193_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y193_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y193_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y193_IOB_X0Y194_IBUF (
.I(LIOB33_X0Y193_IOB_X0Y194_IPAD),
.O(LIOB33_X0Y193_IOB_X0Y194_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y195_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y195_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y195_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y195_IOB_X0Y196_IBUF (
.I(LIOB33_X0Y195_IOB_X0Y196_IPAD),
.O(LIOB33_X0Y195_IOB_X0Y196_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y197_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y197_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y197_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y197_IOB_X0Y198_IBUF (
.I(LIOB33_X0Y197_IOB_X0Y198_IPAD),
.O(LIOB33_X0Y197_IOB_X0Y198_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y201_IOB_X0Y201_IBUF (
.I(LIOB33_X0Y201_IOB_X0Y201_IPAD),
.O(LIOB33_X0Y201_IOB_X0Y201_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y201_IOB_X0Y202_IBUF (
.I(LIOB33_X0Y201_IOB_X0Y202_IPAD),
.O(LIOB33_X0Y201_IOB_X0Y202_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y203_IOB_X0Y203_IBUF (
.I(LIOB33_X0Y203_IOB_X0Y203_IPAD),
.O(LIOB33_X0Y203_IOB_X0Y203_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y99_IOB_X0Y99_OBUF (
.I(CLBLL_R_X71Y131_SLICE_X106Y131_CO6),
.O(LIOB33_SING_X0Y99_IOB_X0Y99_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLM_R_X59Y118_SLICE_X88Y118_AO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_CO6),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y150_IOB_X0Y150_IBUF (
.I(LIOB33_SING_X0Y150_IOB_X0Y150_IPAD),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y199_IOB_X0Y199_IBUF (
.I(LIOB33_SING_X0Y199_IOB_X0Y199_IPAD),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y200_IOB_X0Y200_IBUF (
.I(LIOB33_SING_X0Y200_IOB_X0Y200_IPAD),
.O(LIOB33_SING_X0Y200_IOB_X0Y200_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y51_IOB_X1Y51_IBUF (
.I(RIOB33_X105Y51_IOB_X1Y51_IPAD),
.O(RIOB33_X105Y51_IOB_X1Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y51_IOB_X1Y52_IBUF (
.I(RIOB33_X105Y51_IOB_X1Y52_IPAD),
.O(RIOB33_X105Y51_IOB_X1Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y53_IOB_X1Y53_IBUF (
.I(RIOB33_X105Y53_IOB_X1Y53_IPAD),
.O(RIOB33_X105Y53_IOB_X1Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y53_IOB_X1Y54_IBUF (
.I(RIOB33_X105Y53_IOB_X1Y54_IPAD),
.O(RIOB33_X105Y53_IOB_X1Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y55_IOB_X1Y55_IBUF (
.I(RIOB33_X105Y55_IOB_X1Y55_IPAD),
.O(RIOB33_X105Y55_IOB_X1Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y55_IOB_X1Y56_IBUF (
.I(RIOB33_X105Y55_IOB_X1Y56_IPAD),
.O(RIOB33_X105Y55_IOB_X1Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y57_IOB_X1Y57_IBUF (
.I(RIOB33_X105Y57_IOB_X1Y57_IPAD),
.O(RIOB33_X105Y57_IOB_X1Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y57_IOB_X1Y58_IBUF (
.I(RIOB33_X105Y57_IOB_X1Y58_IPAD),
.O(RIOB33_X105Y57_IOB_X1Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y59_IOB_X1Y59_IBUF (
.I(RIOB33_X105Y59_IOB_X1Y59_IPAD),
.O(RIOB33_X105Y59_IOB_X1Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y59_IOB_X1Y60_IBUF (
.I(RIOB33_X105Y59_IOB_X1Y60_IPAD),
.O(RIOB33_X105Y59_IOB_X1Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y61_IOB_X1Y61_IBUF (
.I(RIOB33_X105Y61_IOB_X1Y61_IPAD),
.O(RIOB33_X105Y61_IOB_X1Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y61_IOB_X1Y62_IBUF (
.I(RIOB33_X105Y61_IOB_X1Y62_IPAD),
.O(RIOB33_X105Y61_IOB_X1Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y63_IOB_X1Y63_IBUF (
.I(RIOB33_X105Y63_IOB_X1Y63_IPAD),
.O(RIOB33_X105Y63_IOB_X1Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y63_IOB_X1Y64_IBUF (
.I(RIOB33_X105Y63_IOB_X1Y64_IPAD),
.O(RIOB33_X105Y63_IOB_X1Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y65_IOB_X1Y65_IBUF (
.I(RIOB33_X105Y65_IOB_X1Y65_IPAD),
.O(RIOB33_X105Y65_IOB_X1Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y65_IOB_X1Y66_IBUF (
.I(RIOB33_X105Y65_IOB_X1Y66_IPAD),
.O(RIOB33_X105Y65_IOB_X1Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y67_IOB_X1Y67_IBUF (
.I(RIOB33_X105Y67_IOB_X1Y67_IPAD),
.O(RIOB33_X105Y67_IOB_X1Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y67_IOB_X1Y68_IBUF (
.I(RIOB33_X105Y67_IOB_X1Y68_IPAD),
.O(RIOB33_X105Y67_IOB_X1Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y69_IOB_X1Y69_IBUF (
.I(RIOB33_X105Y69_IOB_X1Y69_IPAD),
.O(RIOB33_X105Y69_IOB_X1Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y69_IOB_X1Y70_IBUF (
.I(RIOB33_X105Y69_IOB_X1Y70_IPAD),
.O(RIOB33_X105Y69_IOB_X1Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y71_IOB_X1Y71_IBUF (
.I(RIOB33_X105Y71_IOB_X1Y71_IPAD),
.O(RIOB33_X105Y71_IOB_X1Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y71_IOB_X1Y72_IBUF (
.I(RIOB33_X105Y71_IOB_X1Y72_IPAD),
.O(RIOB33_X105Y71_IOB_X1Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y73_IOB_X1Y73_IBUF (
.I(RIOB33_X105Y73_IOB_X1Y73_IPAD),
.O(RIOB33_X105Y73_IOB_X1Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y73_IOB_X1Y74_IBUF (
.I(RIOB33_X105Y73_IOB_X1Y74_IPAD),
.O(RIOB33_X105Y73_IOB_X1Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y75_IOB_X1Y75_IBUF (
.I(RIOB33_X105Y75_IOB_X1Y75_IPAD),
.O(RIOB33_X105Y75_IOB_X1Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y75_IOB_X1Y76_IBUF (
.I(RIOB33_X105Y75_IOB_X1Y76_IPAD),
.O(RIOB33_X105Y75_IOB_X1Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y77_IOB_X1Y77_IBUF (
.I(RIOB33_X105Y77_IOB_X1Y77_IPAD),
.O(RIOB33_X105Y77_IOB_X1Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y77_IOB_X1Y78_IBUF (
.I(RIOB33_X105Y77_IOB_X1Y78_IPAD),
.O(RIOB33_X105Y77_IOB_X1Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y79_IOB_X1Y79_IBUF (
.I(RIOB33_X105Y79_IOB_X1Y79_IPAD),
.O(RIOB33_X105Y79_IOB_X1Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y79_IOB_X1Y80_IBUF (
.I(RIOB33_X105Y79_IOB_X1Y80_IPAD),
.O(RIOB33_X105Y79_IOB_X1Y80_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y81_IOB_X1Y81_IBUF (
.I(RIOB33_X105Y81_IOB_X1Y81_IPAD),
.O(RIOB33_X105Y81_IOB_X1Y81_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y81_IOB_X1Y82_IBUF (
.I(RIOB33_X105Y81_IOB_X1Y82_IPAD),
.O(RIOB33_X105Y81_IOB_X1Y82_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y83_IOB_X1Y83_IBUF (
.I(RIOB33_X105Y83_IOB_X1Y83_IPAD),
.O(RIOB33_X105Y83_IOB_X1Y83_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y83_IOB_X1Y84_IBUF (
.I(RIOB33_X105Y83_IOB_X1Y84_IPAD),
.O(RIOB33_X105Y83_IOB_X1Y84_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y85_IOB_X1Y85_IBUF (
.I(RIOB33_X105Y85_IOB_X1Y85_IPAD),
.O(RIOB33_X105Y85_IOB_X1Y85_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y85_IOB_X1Y86_IBUF (
.I(RIOB33_X105Y85_IOB_X1Y86_IPAD),
.O(RIOB33_X105Y85_IOB_X1Y86_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y87_IOB_X1Y87_IBUF (
.I(RIOB33_X105Y87_IOB_X1Y87_IPAD),
.O(RIOB33_X105Y87_IOB_X1Y87_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y87_IOB_X1Y88_IBUF (
.I(RIOB33_X105Y87_IOB_X1Y88_IPAD),
.O(RIOB33_X105Y87_IOB_X1Y88_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y89_IOB_X1Y89_IBUF (
.I(RIOB33_X105Y89_IOB_X1Y89_IPAD),
.O(RIOB33_X105Y89_IOB_X1Y89_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y89_IOB_X1Y90_IBUF (
.I(RIOB33_X105Y89_IOB_X1Y90_IPAD),
.O(RIOB33_X105Y89_IOB_X1Y90_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y91_IOB_X1Y91_IBUF (
.I(RIOB33_X105Y91_IOB_X1Y91_IPAD),
.O(RIOB33_X105Y91_IOB_X1Y91_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y91_IOB_X1Y92_IBUF (
.I(RIOB33_X105Y91_IOB_X1Y92_IPAD),
.O(RIOB33_X105Y91_IOB_X1Y92_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y93_IOB_X1Y93_IBUF (
.I(RIOB33_X105Y93_IOB_X1Y93_IPAD),
.O(RIOB33_X105Y93_IOB_X1Y93_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y93_IOB_X1Y94_IBUF (
.I(RIOB33_X105Y93_IOB_X1Y94_IPAD),
.O(RIOB33_X105Y93_IOB_X1Y94_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y95_IOB_X1Y95_IBUF (
.I(RIOB33_X105Y95_IOB_X1Y95_IPAD),
.O(RIOB33_X105Y95_IOB_X1Y95_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y95_IOB_X1Y96_IBUF (
.I(RIOB33_X105Y95_IOB_X1Y96_IPAD),
.O(RIOB33_X105Y95_IOB_X1Y96_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y97_IOB_X1Y97_IBUF (
.I(RIOB33_X105Y97_IOB_X1Y97_IPAD),
.O(RIOB33_X105Y97_IOB_X1Y97_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y97_IOB_X1Y98_IBUF (
.I(RIOB33_X105Y97_IOB_X1Y98_IPAD),
.O(RIOB33_X105Y97_IOB_X1Y98_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y151_IOB_X1Y151_IBUF (
.I(RIOB33_X105Y151_IOB_X1Y151_IPAD),
.O(RIOB33_X105Y151_IOB_X1Y151_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y151_IOB_X1Y152_IBUF (
.I(RIOB33_X105Y151_IOB_X1Y152_IPAD),
.O(RIOB33_X105Y151_IOB_X1Y152_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y153_IOB_X1Y153_IBUF (
.I(RIOB33_X105Y153_IOB_X1Y153_IPAD),
.O(RIOB33_X105Y153_IOB_X1Y153_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y153_IOB_X1Y154_IBUF (
.I(RIOB33_X105Y153_IOB_X1Y154_IPAD),
.O(RIOB33_X105Y153_IOB_X1Y154_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y155_IOB_X1Y155_IBUF (
.I(RIOB33_X105Y155_IOB_X1Y155_IPAD),
.O(RIOB33_X105Y155_IOB_X1Y155_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y155_IOB_X1Y156_IBUF (
.I(RIOB33_X105Y155_IOB_X1Y156_IPAD),
.O(RIOB33_X105Y155_IOB_X1Y156_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y157_IOB_X1Y157_IBUF (
.I(RIOB33_X105Y157_IOB_X1Y157_IPAD),
.O(RIOB33_X105Y157_IOB_X1Y157_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y157_IOB_X1Y158_IBUF (
.I(RIOB33_X105Y157_IOB_X1Y158_IPAD),
.O(RIOB33_X105Y157_IOB_X1Y158_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y159_IOB_X1Y159_IBUF (
.I(RIOB33_X105Y159_IOB_X1Y159_IPAD),
.O(RIOB33_X105Y159_IOB_X1Y159_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y159_IOB_X1Y160_IBUF (
.I(RIOB33_X105Y159_IOB_X1Y160_IPAD),
.O(RIOB33_X105Y159_IOB_X1Y160_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y161_IOB_X1Y161_IBUF (
.I(RIOB33_X105Y161_IOB_X1Y161_IPAD),
.O(RIOB33_X105Y161_IOB_X1Y161_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y161_IOB_X1Y162_IBUF (
.I(RIOB33_X105Y161_IOB_X1Y162_IPAD),
.O(RIOB33_X105Y161_IOB_X1Y162_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y163_IOB_X1Y163_IBUF (
.I(RIOB33_X105Y163_IOB_X1Y163_IPAD),
.O(RIOB33_X105Y163_IOB_X1Y163_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y163_IOB_X1Y164_IBUF (
.I(RIOB33_X105Y163_IOB_X1Y164_IPAD),
.O(RIOB33_X105Y163_IOB_X1Y164_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y165_IOB_X1Y165_IBUF (
.I(RIOB33_X105Y165_IOB_X1Y165_IPAD),
.O(RIOB33_X105Y165_IOB_X1Y165_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y165_IOB_X1Y166_IBUF (
.I(RIOB33_X105Y165_IOB_X1Y166_IPAD),
.O(RIOB33_X105Y165_IOB_X1Y166_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y167_IOB_X1Y167_IBUF (
.I(RIOB33_X105Y167_IOB_X1Y167_IPAD),
.O(RIOB33_X105Y167_IOB_X1Y167_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y167_IOB_X1Y168_IBUF (
.I(RIOB33_X105Y167_IOB_X1Y168_IPAD),
.O(RIOB33_X105Y167_IOB_X1Y168_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y169_IOB_X1Y169_IBUF (
.I(RIOB33_X105Y169_IOB_X1Y169_IPAD),
.O(RIOB33_X105Y169_IOB_X1Y169_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y169_IOB_X1Y170_IBUF (
.I(RIOB33_X105Y169_IOB_X1Y170_IPAD),
.O(RIOB33_X105Y169_IOB_X1Y170_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y171_IOB_X1Y171_IBUF (
.I(RIOB33_X105Y171_IOB_X1Y171_IPAD),
.O(RIOB33_X105Y171_IOB_X1Y171_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y171_IOB_X1Y172_IBUF (
.I(RIOB33_X105Y171_IOB_X1Y172_IPAD),
.O(RIOB33_X105Y171_IOB_X1Y172_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y173_IOB_X1Y173_IBUF (
.I(RIOB33_X105Y173_IOB_X1Y173_IPAD),
.O(RIOB33_X105Y173_IOB_X1Y173_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y173_IOB_X1Y174_IBUF (
.I(RIOB33_X105Y173_IOB_X1Y174_IPAD),
.O(RIOB33_X105Y173_IOB_X1Y174_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y175_IOB_X1Y175_IBUF (
.I(RIOB33_X105Y175_IOB_X1Y175_IPAD),
.O(RIOB33_X105Y175_IOB_X1Y175_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y175_IOB_X1Y176_IBUF (
.I(RIOB33_X105Y175_IOB_X1Y176_IPAD),
.O(RIOB33_X105Y175_IOB_X1Y176_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y177_IOB_X1Y177_IBUF (
.I(RIOB33_X105Y177_IOB_X1Y177_IPAD),
.O(RIOB33_X105Y177_IOB_X1Y177_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y177_IOB_X1Y178_IBUF (
.I(RIOB33_X105Y177_IOB_X1Y178_IPAD),
.O(RIOB33_X105Y177_IOB_X1Y178_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y179_IOB_X1Y179_IBUF (
.I(RIOB33_X105Y179_IOB_X1Y179_IPAD),
.O(RIOB33_X105Y179_IOB_X1Y179_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y179_IOB_X1Y180_IBUF (
.I(RIOB33_X105Y179_IOB_X1Y180_IPAD),
.O(RIOB33_X105Y179_IOB_X1Y180_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y181_IOB_X1Y181_IBUF (
.I(RIOB33_X105Y181_IOB_X1Y181_IPAD),
.O(RIOB33_X105Y181_IOB_X1Y181_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y181_IOB_X1Y182_IBUF (
.I(RIOB33_X105Y181_IOB_X1Y182_IPAD),
.O(RIOB33_X105Y181_IOB_X1Y182_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y183_IOB_X1Y183_IBUF (
.I(RIOB33_X105Y183_IOB_X1Y183_IPAD),
.O(RIOB33_X105Y183_IOB_X1Y183_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y183_IOB_X1Y184_IBUF (
.I(RIOB33_X105Y183_IOB_X1Y184_IPAD),
.O(RIOB33_X105Y183_IOB_X1Y184_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y185_IOB_X1Y185_IBUF (
.I(RIOB33_X105Y185_IOB_X1Y185_IPAD),
.O(RIOB33_X105Y185_IOB_X1Y185_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y185_IOB_X1Y186_IBUF (
.I(RIOB33_X105Y185_IOB_X1Y186_IPAD),
.O(RIOB33_X105Y185_IOB_X1Y186_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y187_IOB_X1Y187_IBUF (
.I(RIOB33_X105Y187_IOB_X1Y187_IPAD),
.O(RIOB33_X105Y187_IOB_X1Y187_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y187_IOB_X1Y188_IBUF (
.I(RIOB33_X105Y187_IOB_X1Y188_IPAD),
.O(RIOB33_X105Y187_IOB_X1Y188_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y189_IOB_X1Y189_IBUF (
.I(RIOB33_X105Y189_IOB_X1Y189_IPAD),
.O(RIOB33_X105Y189_IOB_X1Y189_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y189_IOB_X1Y190_IBUF (
.I(RIOB33_X105Y189_IOB_X1Y190_IPAD),
.O(RIOB33_X105Y189_IOB_X1Y190_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y191_IOB_X1Y191_IBUF (
.I(RIOB33_X105Y191_IOB_X1Y191_IPAD),
.O(RIOB33_X105Y191_IOB_X1Y191_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y191_IOB_X1Y192_IBUF (
.I(RIOB33_X105Y191_IOB_X1Y192_IPAD),
.O(RIOB33_X105Y191_IOB_X1Y192_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y193_IOB_X1Y193_IBUF (
.I(RIOB33_X105Y193_IOB_X1Y193_IPAD),
.O(RIOB33_X105Y193_IOB_X1Y193_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y193_IOB_X1Y194_IBUF (
.I(RIOB33_X105Y193_IOB_X1Y194_IPAD),
.O(RIOB33_X105Y193_IOB_X1Y194_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y195_IOB_X1Y195_IBUF (
.I(RIOB33_X105Y195_IOB_X1Y195_IPAD),
.O(RIOB33_X105Y195_IOB_X1Y195_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y195_IOB_X1Y196_IBUF (
.I(RIOB33_X105Y195_IOB_X1Y196_IPAD),
.O(RIOB33_X105Y195_IOB_X1Y196_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y197_IOB_X1Y197_IBUF (
.I(RIOB33_X105Y197_IOB_X1Y197_IPAD),
.O(RIOB33_X105Y197_IOB_X1Y197_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y197_IOB_X1Y198_IBUF (
.I(RIOB33_X105Y197_IOB_X1Y198_IPAD),
.O(RIOB33_X105Y197_IOB_X1Y198_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y50_IOB_X1Y50_IBUF (
.I(RIOB33_SING_X105Y50_IOB_X1Y50_IPAD),
.O(RIOB33_SING_X105Y50_IOB_X1Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y99_IOB_X1Y99_IBUF (
.I(RIOB33_SING_X105Y99_IOB_X1Y99_IPAD),
.O(RIOB33_SING_X105Y99_IOB_X1Y99_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y150_IOB_X1Y150_IBUF (
.I(RIOB33_SING_X105Y150_IOB_X1Y150_IPAD),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y199_IOB_X1Y199_IBUF (
.I(RIOB33_SING_X105Y199_IOB_X1Y199_IPAD),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_I)
  );
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_BMUX = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_AMUX = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C = CLBLL_L_X2Y123_SLICE_X1Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D = CLBLL_L_X2Y123_SLICE_X1Y123_DO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B = CLBLL_L_X2Y124_SLICE_X0Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_DMUX = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B = CLBLL_L_X2Y124_SLICE_X1Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_A = CLBLL_R_X71Y116_SLICE_X106Y116_AO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_B = CLBLL_R_X71Y116_SLICE_X106Y116_BO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_C = CLBLL_R_X71Y116_SLICE_X106Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_D = CLBLL_R_X71Y116_SLICE_X106Y116_DO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_BMUX = CLBLL_R_X71Y116_SLICE_X106Y116_F8MUX_O;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_A = CLBLL_R_X71Y116_SLICE_X107Y116_AO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_B = CLBLL_R_X71Y116_SLICE_X107Y116_BO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_C = CLBLL_R_X71Y116_SLICE_X107Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_D = CLBLL_R_X71Y116_SLICE_X107Y116_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A = CLBLL_R_X71Y117_SLICE_X106Y117_AO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B = CLBLL_R_X71Y117_SLICE_X106Y117_BO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C = CLBLL_R_X71Y117_SLICE_X106Y117_CO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D = CLBLL_R_X71Y117_SLICE_X106Y117_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_AMUX = CLBLL_R_X71Y117_SLICE_X106Y117_F7AMUX_O;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_CMUX = CLBLL_R_X71Y117_SLICE_X106Y117_F7BMUX_O;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A = CLBLL_R_X71Y117_SLICE_X107Y117_AO6;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B = CLBLL_R_X71Y117_SLICE_X107Y117_BO6;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C = CLBLL_R_X71Y117_SLICE_X107Y117_CO6;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D = CLBLL_R_X71Y117_SLICE_X107Y117_DO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_A = CLBLL_R_X71Y118_SLICE_X106Y118_AO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_B = CLBLL_R_X71Y118_SLICE_X106Y118_BO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_C = CLBLL_R_X71Y118_SLICE_X106Y118_CO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_D = CLBLL_R_X71Y118_SLICE_X106Y118_DO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_A = CLBLL_R_X71Y118_SLICE_X107Y118_AO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_B = CLBLL_R_X71Y118_SLICE_X107Y118_BO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_C = CLBLL_R_X71Y118_SLICE_X107Y118_CO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_D = CLBLL_R_X71Y118_SLICE_X107Y118_DO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_BMUX = CLBLL_R_X71Y118_SLICE_X107Y118_F8MUX_O;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A = CLBLL_R_X71Y119_SLICE_X106Y119_AO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B = CLBLL_R_X71Y119_SLICE_X106Y119_BO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C = CLBLL_R_X71Y119_SLICE_X106Y119_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D = CLBLL_R_X71Y119_SLICE_X106Y119_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A = CLBLL_R_X71Y119_SLICE_X107Y119_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B = CLBLL_R_X71Y119_SLICE_X107Y119_BO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C = CLBLL_R_X71Y119_SLICE_X107Y119_CO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D = CLBLL_R_X71Y119_SLICE_X107Y119_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_AMUX = CLBLL_R_X71Y119_SLICE_X107Y119_F7AMUX_O;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_CMUX = CLBLL_R_X71Y119_SLICE_X107Y119_F7BMUX_O;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_A = CLBLL_R_X71Y120_SLICE_X106Y120_AO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_B = CLBLL_R_X71Y120_SLICE_X106Y120_BO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_C = CLBLL_R_X71Y120_SLICE_X106Y120_CO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_D = CLBLL_R_X71Y120_SLICE_X106Y120_DO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_AMUX = CLBLL_R_X71Y120_SLICE_X106Y120_F7AMUX_O;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_CMUX = CLBLL_R_X71Y120_SLICE_X106Y120_F7BMUX_O;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_A = CLBLL_R_X71Y120_SLICE_X107Y120_AO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_B = CLBLL_R_X71Y120_SLICE_X107Y120_BO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_C = CLBLL_R_X71Y120_SLICE_X107Y120_CO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_D = CLBLL_R_X71Y120_SLICE_X107Y120_DO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A = CLBLL_R_X71Y121_SLICE_X106Y121_AO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B = CLBLL_R_X71Y121_SLICE_X106Y121_BO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C = CLBLL_R_X71Y121_SLICE_X106Y121_CO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D = CLBLL_R_X71Y121_SLICE_X106Y121_DO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_AMUX = CLBLL_R_X71Y121_SLICE_X106Y121_F7AMUX_O;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_CMUX = CLBLL_R_X71Y121_SLICE_X106Y121_F7BMUX_O;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A = CLBLL_R_X71Y121_SLICE_X107Y121_AO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B = CLBLL_R_X71Y121_SLICE_X107Y121_BO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C = CLBLL_R_X71Y121_SLICE_X107Y121_CO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D = CLBLL_R_X71Y121_SLICE_X107Y121_DO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_BMUX = CLBLL_R_X71Y121_SLICE_X107Y121_F8MUX_O;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_A = CLBLL_R_X71Y122_SLICE_X106Y122_AO6;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_B = CLBLL_R_X71Y122_SLICE_X106Y122_BO6;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_C = CLBLL_R_X71Y122_SLICE_X106Y122_CO6;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_D = CLBLL_R_X71Y122_SLICE_X106Y122_DO6;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_AMUX = CLBLL_R_X71Y122_SLICE_X106Y122_AO6;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_A = CLBLL_R_X71Y122_SLICE_X107Y122_AO6;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_B = CLBLL_R_X71Y122_SLICE_X107Y122_BO6;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_C = CLBLL_R_X71Y122_SLICE_X107Y122_CO6;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_D = CLBLL_R_X71Y122_SLICE_X107Y122_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A = CLBLL_R_X71Y125_SLICE_X106Y125_AO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B = CLBLL_R_X71Y125_SLICE_X106Y125_BO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C = CLBLL_R_X71Y125_SLICE_X106Y125_CO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D = CLBLL_R_X71Y125_SLICE_X106Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A = CLBLL_R_X71Y125_SLICE_X107Y125_AO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B = CLBLL_R_X71Y125_SLICE_X107Y125_BO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D = CLBLL_R_X71Y125_SLICE_X107Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_AMUX = CLBLL_R_X71Y125_SLICE_X107Y125_F7AMUX_O;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A = CLBLL_R_X71Y126_SLICE_X106Y126_AO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B = CLBLL_R_X71Y126_SLICE_X106Y126_BO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C = CLBLL_R_X71Y126_SLICE_X106Y126_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D = CLBLL_R_X71Y126_SLICE_X106Y126_DO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A = CLBLL_R_X71Y126_SLICE_X107Y126_AO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B = CLBLL_R_X71Y126_SLICE_X107Y126_BO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C = CLBLL_R_X71Y126_SLICE_X107Y126_CO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D = CLBLL_R_X71Y126_SLICE_X107Y126_DO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_AMUX = CLBLL_R_X71Y126_SLICE_X107Y126_F7AMUX_O;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A = CLBLL_R_X71Y127_SLICE_X106Y127_AO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B = CLBLL_R_X71Y127_SLICE_X106Y127_BO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C = CLBLL_R_X71Y127_SLICE_X106Y127_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D = CLBLL_R_X71Y127_SLICE_X106Y127_DO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A = CLBLL_R_X71Y127_SLICE_X107Y127_AO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B = CLBLL_R_X71Y127_SLICE_X107Y127_BO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C = CLBLL_R_X71Y127_SLICE_X107Y127_CO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D = CLBLL_R_X71Y127_SLICE_X107Y127_DO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A = CLBLL_R_X71Y128_SLICE_X106Y128_AO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B = CLBLL_R_X71Y128_SLICE_X106Y128_BO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D = CLBLL_R_X71Y128_SLICE_X106Y128_DO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_AMUX = CLBLL_R_X71Y128_SLICE_X106Y128_AO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_CMUX = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A = CLBLL_R_X71Y128_SLICE_X107Y128_AO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B = CLBLL_R_X71Y128_SLICE_X107Y128_BO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C = CLBLL_R_X71Y128_SLICE_X107Y128_CO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D = CLBLL_R_X71Y128_SLICE_X107Y128_DO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A = CLBLL_R_X71Y129_SLICE_X106Y129_AO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B = CLBLL_R_X71Y129_SLICE_X106Y129_BO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C = CLBLL_R_X71Y129_SLICE_X106Y129_CO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D = CLBLL_R_X71Y129_SLICE_X106Y129_DO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A = CLBLL_R_X71Y129_SLICE_X107Y129_AO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B = CLBLL_R_X71Y129_SLICE_X107Y129_BO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C = CLBLL_R_X71Y129_SLICE_X107Y129_CO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D = CLBLL_R_X71Y129_SLICE_X107Y129_DO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A = CLBLL_R_X71Y131_SLICE_X106Y131_AO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B = CLBLL_R_X71Y131_SLICE_X106Y131_BO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C = CLBLL_R_X71Y131_SLICE_X106Y131_CO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D = CLBLL_R_X71Y131_SLICE_X106Y131_DO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A = CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B = CLBLL_R_X71Y131_SLICE_X107Y131_BO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C = CLBLL_R_X71Y131_SLICE_X107Y131_CO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D = CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_AMUX = CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_CMUX = CLBLL_R_X71Y131_SLICE_X107Y131_CO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_A = CLBLL_R_X73Y114_SLICE_X110Y114_AO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_B = CLBLL_R_X73Y114_SLICE_X110Y114_BO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_C = CLBLL_R_X73Y114_SLICE_X110Y114_CO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_D = CLBLL_R_X73Y114_SLICE_X110Y114_DO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_BMUX = CLBLL_R_X73Y114_SLICE_X110Y114_F8MUX_O;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_A = CLBLL_R_X73Y114_SLICE_X111Y114_AO6;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_B = CLBLL_R_X73Y114_SLICE_X111Y114_BO6;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_C = CLBLL_R_X73Y114_SLICE_X111Y114_CO6;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_D = CLBLL_R_X73Y114_SLICE_X111Y114_DO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_A = CLBLL_R_X73Y115_SLICE_X110Y115_AO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_B = CLBLL_R_X73Y115_SLICE_X110Y115_BO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_C = CLBLL_R_X73Y115_SLICE_X110Y115_CO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_D = CLBLL_R_X73Y115_SLICE_X110Y115_DO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_AMUX = CLBLL_R_X73Y115_SLICE_X110Y115_F7AMUX_O;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_A = CLBLL_R_X73Y115_SLICE_X111Y115_AO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_B = CLBLL_R_X73Y115_SLICE_X111Y115_BO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_C = CLBLL_R_X73Y115_SLICE_X111Y115_CO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_D = CLBLL_R_X73Y115_SLICE_X111Y115_DO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_BMUX = CLBLL_R_X73Y115_SLICE_X111Y115_F8MUX_O;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_A = CLBLL_R_X73Y116_SLICE_X110Y116_AO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_B = CLBLL_R_X73Y116_SLICE_X110Y116_BO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_C = CLBLL_R_X73Y116_SLICE_X110Y116_CO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_D = CLBLL_R_X73Y116_SLICE_X110Y116_DO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_AMUX = CLBLL_R_X73Y116_SLICE_X110Y116_F7AMUX_O;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_A = CLBLL_R_X73Y116_SLICE_X111Y116_AO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_B = CLBLL_R_X73Y116_SLICE_X111Y116_BO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_C = CLBLL_R_X73Y116_SLICE_X111Y116_CO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_D = CLBLL_R_X73Y116_SLICE_X111Y116_DO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_BMUX = CLBLL_R_X73Y116_SLICE_X111Y116_F8MUX_O;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A = CLBLL_R_X73Y118_SLICE_X110Y118_AO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B = CLBLL_R_X73Y118_SLICE_X110Y118_BO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C = CLBLL_R_X73Y118_SLICE_X110Y118_CO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D = CLBLL_R_X73Y118_SLICE_X110Y118_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_BMUX = CLBLL_R_X73Y118_SLICE_X110Y118_F8MUX_O;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A = CLBLL_R_X73Y118_SLICE_X111Y118_AO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B = CLBLL_R_X73Y118_SLICE_X111Y118_BO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C = CLBLL_R_X73Y118_SLICE_X111Y118_CO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D = CLBLL_R_X73Y118_SLICE_X111Y118_DO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_AMUX = CLBLL_R_X73Y118_SLICE_X111Y118_F7AMUX_O;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A = CLBLL_R_X73Y119_SLICE_X110Y119_AO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B = CLBLL_R_X73Y119_SLICE_X110Y119_BO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C = CLBLL_R_X73Y119_SLICE_X110Y119_CO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D = CLBLL_R_X73Y119_SLICE_X110Y119_DO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_BMUX = CLBLL_R_X73Y119_SLICE_X110Y119_F8MUX_O;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A = CLBLL_R_X73Y119_SLICE_X111Y119_AO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B = CLBLL_R_X73Y119_SLICE_X111Y119_BO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C = CLBLL_R_X73Y119_SLICE_X111Y119_CO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_AMUX = CLBLL_R_X73Y119_SLICE_X111Y119_F7AMUX_O;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_A = CLBLL_R_X73Y120_SLICE_X110Y120_AO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_B = CLBLL_R_X73Y120_SLICE_X110Y120_BO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_C = CLBLL_R_X73Y120_SLICE_X110Y120_CO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_D = CLBLL_R_X73Y120_SLICE_X110Y120_DO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_AMUX = CLBLL_R_X73Y120_SLICE_X110Y120_F7AMUX_O;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_CMUX = CLBLL_R_X73Y120_SLICE_X110Y120_F7BMUX_O;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_A = CLBLL_R_X73Y120_SLICE_X111Y120_AO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_B = CLBLL_R_X73Y120_SLICE_X111Y120_BO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_C = CLBLL_R_X73Y120_SLICE_X111Y120_CO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_D = CLBLL_R_X73Y120_SLICE_X111Y120_DO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_AMUX = CLBLL_R_X73Y120_SLICE_X111Y120_F7AMUX_O;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A = CLBLL_R_X73Y121_SLICE_X110Y121_AO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B = CLBLL_R_X73Y121_SLICE_X110Y121_BO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C = CLBLL_R_X73Y121_SLICE_X110Y121_CO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D = CLBLL_R_X73Y121_SLICE_X110Y121_DO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_AMUX = CLBLL_R_X73Y121_SLICE_X110Y121_F7AMUX_O;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A = CLBLL_R_X73Y121_SLICE_X111Y121_AO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B = CLBLL_R_X73Y121_SLICE_X111Y121_BO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C = CLBLL_R_X73Y121_SLICE_X111Y121_CO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D = CLBLL_R_X73Y121_SLICE_X111Y121_DO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_AMUX = CLBLL_R_X73Y121_SLICE_X111Y121_F7AMUX_O;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_CMUX = CLBLL_R_X73Y121_SLICE_X111Y121_F7BMUX_O;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A = CLBLL_R_X73Y122_SLICE_X110Y122_AO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B = CLBLL_R_X73Y122_SLICE_X110Y122_BO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C = CLBLL_R_X73Y122_SLICE_X110Y122_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D = CLBLL_R_X73Y122_SLICE_X110Y122_DO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A = CLBLL_R_X73Y122_SLICE_X111Y122_AO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B = CLBLL_R_X73Y122_SLICE_X111Y122_BO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C = CLBLL_R_X73Y122_SLICE_X111Y122_CO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D = CLBLL_R_X73Y122_SLICE_X111Y122_DO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A = CLBLL_R_X73Y123_SLICE_X110Y123_AO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B = CLBLL_R_X73Y123_SLICE_X110Y123_BO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C = CLBLL_R_X73Y123_SLICE_X110Y123_CO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D = CLBLL_R_X73Y123_SLICE_X110Y123_DO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_AMUX = CLBLL_R_X73Y123_SLICE_X110Y123_F7AMUX_O;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A = CLBLL_R_X73Y123_SLICE_X111Y123_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B = CLBLL_R_X73Y123_SLICE_X111Y123_BO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C = CLBLL_R_X73Y123_SLICE_X111Y123_CO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D = CLBLL_R_X73Y123_SLICE_X111Y123_DO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_BMUX = CLBLL_R_X73Y123_SLICE_X111Y123_F8MUX_O;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A = CLBLL_R_X73Y124_SLICE_X110Y124_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B = CLBLL_R_X73Y124_SLICE_X110Y124_BO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C = CLBLL_R_X73Y124_SLICE_X110Y124_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D = CLBLL_R_X73Y124_SLICE_X110Y124_DO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_BMUX = CLBLL_R_X73Y124_SLICE_X110Y124_F8MUX_O;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A = CLBLL_R_X73Y124_SLICE_X111Y124_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B = CLBLL_R_X73Y124_SLICE_X111Y124_BO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C = CLBLL_R_X73Y124_SLICE_X111Y124_CO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D = CLBLL_R_X73Y124_SLICE_X111Y124_DO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_AMUX = CLBLL_R_X73Y124_SLICE_X111Y124_F7AMUX_O;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_CMUX = CLBLL_R_X73Y124_SLICE_X111Y124_F7BMUX_O;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A = CLBLL_R_X73Y125_SLICE_X110Y125_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B = CLBLL_R_X73Y125_SLICE_X110Y125_BO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C = CLBLL_R_X73Y125_SLICE_X110Y125_CO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D = CLBLL_R_X73Y125_SLICE_X110Y125_DO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_BMUX = CLBLL_R_X73Y125_SLICE_X110Y125_F8MUX_O;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A = CLBLL_R_X73Y125_SLICE_X111Y125_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B = CLBLL_R_X73Y125_SLICE_X111Y125_BO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C = CLBLL_R_X73Y125_SLICE_X111Y125_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D = CLBLL_R_X73Y125_SLICE_X111Y125_DO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_BMUX = CLBLL_R_X73Y125_SLICE_X111Y125_F8MUX_O;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A = CLBLL_R_X73Y126_SLICE_X110Y126_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B = CLBLL_R_X73Y126_SLICE_X110Y126_BO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C = CLBLL_R_X73Y126_SLICE_X110Y126_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D = CLBLL_R_X73Y126_SLICE_X110Y126_DO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_BMUX = CLBLL_R_X73Y126_SLICE_X110Y126_F8MUX_O;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A = CLBLL_R_X73Y126_SLICE_X111Y126_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B = CLBLL_R_X73Y126_SLICE_X111Y126_BO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C = CLBLL_R_X73Y126_SLICE_X111Y126_CO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D = CLBLL_R_X73Y126_SLICE_X111Y126_DO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_AMUX = CLBLL_R_X73Y126_SLICE_X111Y126_F7AMUX_O;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_CMUX = CLBLL_R_X73Y126_SLICE_X111Y126_F7BMUX_O;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A = CLBLL_R_X73Y127_SLICE_X110Y127_AO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B = CLBLL_R_X73Y127_SLICE_X110Y127_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C = CLBLL_R_X73Y127_SLICE_X110Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D = CLBLL_R_X73Y127_SLICE_X110Y127_DO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_BMUX = CLBLL_R_X73Y127_SLICE_X110Y127_F8MUX_O;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A = CLBLL_R_X73Y127_SLICE_X111Y127_AO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B = CLBLL_R_X73Y127_SLICE_X111Y127_BO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C = CLBLL_R_X73Y127_SLICE_X111Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D = CLBLL_R_X73Y127_SLICE_X111Y127_DO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_AMUX = CLBLL_R_X73Y127_SLICE_X111Y127_F7AMUX_O;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A = CLBLL_R_X73Y128_SLICE_X110Y128_AO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B = CLBLL_R_X73Y128_SLICE_X110Y128_BO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C = CLBLL_R_X73Y128_SLICE_X110Y128_CO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D = CLBLL_R_X73Y128_SLICE_X110Y128_DO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_BMUX = CLBLL_R_X73Y128_SLICE_X110Y128_F8MUX_O;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A = CLBLL_R_X73Y128_SLICE_X111Y128_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B = CLBLL_R_X73Y128_SLICE_X111Y128_BO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C = CLBLL_R_X73Y128_SLICE_X111Y128_CO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D = CLBLL_R_X73Y128_SLICE_X111Y128_DO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_AMUX = CLBLL_R_X73Y128_SLICE_X111Y128_F7AMUX_O;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_CMUX = CLBLL_R_X73Y128_SLICE_X111Y128_F7BMUX_O;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_A = CLBLL_R_X73Y129_SLICE_X110Y129_AO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_B = CLBLL_R_X73Y129_SLICE_X110Y129_BO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_C = CLBLL_R_X73Y129_SLICE_X110Y129_CO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_D = CLBLL_R_X73Y129_SLICE_X110Y129_DO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_AMUX = CLBLL_R_X73Y129_SLICE_X110Y129_F7AMUX_O;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_A = CLBLL_R_X73Y129_SLICE_X111Y129_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_B = CLBLL_R_X73Y129_SLICE_X111Y129_BO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_C = CLBLL_R_X73Y129_SLICE_X111Y129_CO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_D = CLBLL_R_X73Y129_SLICE_X111Y129_DO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_BMUX = CLBLL_R_X73Y129_SLICE_X111Y129_F8MUX_O;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_A = CLBLL_R_X75Y115_SLICE_X114Y115_AO6;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_B = CLBLL_R_X75Y115_SLICE_X114Y115_BO6;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_C = CLBLL_R_X75Y115_SLICE_X114Y115_CO6;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_D = CLBLL_R_X75Y115_SLICE_X114Y115_DO6;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_AMUX = CLBLL_R_X75Y115_SLICE_X114Y115_F7AMUX_O;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_A = CLBLL_R_X75Y115_SLICE_X115Y115_AO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_B = CLBLL_R_X75Y115_SLICE_X115Y115_BO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_C = CLBLL_R_X75Y115_SLICE_X115Y115_CO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_D = CLBLL_R_X75Y115_SLICE_X115Y115_DO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_BMUX = CLBLL_R_X75Y115_SLICE_X115Y115_F8MUX_O;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_A = CLBLL_R_X75Y116_SLICE_X114Y116_AO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_B = CLBLL_R_X75Y116_SLICE_X114Y116_BO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_C = CLBLL_R_X75Y116_SLICE_X114Y116_CO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_D = CLBLL_R_X75Y116_SLICE_X114Y116_DO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_AMUX = CLBLL_R_X75Y116_SLICE_X114Y116_F7AMUX_O;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_A = CLBLL_R_X75Y116_SLICE_X115Y116_AO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_B = CLBLL_R_X75Y116_SLICE_X115Y116_BO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_C = CLBLL_R_X75Y116_SLICE_X115Y116_CO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_D = CLBLL_R_X75Y116_SLICE_X115Y116_DO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_AMUX = CLBLL_R_X75Y116_SLICE_X115Y116_F7AMUX_O;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_A = CLBLL_R_X75Y117_SLICE_X114Y117_AO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_B = CLBLL_R_X75Y117_SLICE_X114Y117_BO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_C = CLBLL_R_X75Y117_SLICE_X114Y117_CO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_D = CLBLL_R_X75Y117_SLICE_X114Y117_DO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_AMUX = CLBLL_R_X75Y117_SLICE_X114Y117_F7AMUX_O;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_CMUX = CLBLL_R_X75Y117_SLICE_X114Y117_F7BMUX_O;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_A = CLBLL_R_X75Y117_SLICE_X115Y117_AO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_B = CLBLL_R_X75Y117_SLICE_X115Y117_BO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_C = CLBLL_R_X75Y117_SLICE_X115Y117_CO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_D = CLBLL_R_X75Y117_SLICE_X115Y117_DO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_BMUX = CLBLL_R_X75Y117_SLICE_X115Y117_F8MUX_O;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_A = CLBLL_R_X75Y118_SLICE_X114Y118_AO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_B = CLBLL_R_X75Y118_SLICE_X114Y118_BO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_C = CLBLL_R_X75Y118_SLICE_X114Y118_CO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_D = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_AMUX = CLBLL_R_X75Y118_SLICE_X114Y118_F7AMUX_O;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_A = CLBLL_R_X75Y118_SLICE_X115Y118_AO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_B = CLBLL_R_X75Y118_SLICE_X115Y118_BO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_C = CLBLL_R_X75Y118_SLICE_X115Y118_CO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_D = CLBLL_R_X75Y118_SLICE_X115Y118_DO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_BMUX = CLBLL_R_X75Y118_SLICE_X115Y118_F8MUX_O;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_A = CLBLL_R_X75Y119_SLICE_X114Y119_AO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_B = CLBLL_R_X75Y119_SLICE_X114Y119_BO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_C = CLBLL_R_X75Y119_SLICE_X114Y119_CO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_D = CLBLL_R_X75Y119_SLICE_X114Y119_DO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_AMUX = CLBLL_R_X75Y119_SLICE_X114Y119_F7AMUX_O;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_A = CLBLL_R_X75Y119_SLICE_X115Y119_AO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_B = CLBLL_R_X75Y119_SLICE_X115Y119_BO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_C = CLBLL_R_X75Y119_SLICE_X115Y119_CO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_D = CLBLL_R_X75Y119_SLICE_X115Y119_DO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_AMUX = CLBLL_R_X75Y119_SLICE_X115Y119_F7AMUX_O;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_A = CLBLL_R_X75Y120_SLICE_X114Y120_AO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_B = CLBLL_R_X75Y120_SLICE_X114Y120_BO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_C = CLBLL_R_X75Y120_SLICE_X114Y120_CO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_D = CLBLL_R_X75Y120_SLICE_X114Y120_DO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_BMUX = CLBLL_R_X75Y120_SLICE_X114Y120_F8MUX_O;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_A = CLBLL_R_X75Y120_SLICE_X115Y120_AO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_B = CLBLL_R_X75Y120_SLICE_X115Y120_BO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_C = CLBLL_R_X75Y120_SLICE_X115Y120_CO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_D = CLBLL_R_X75Y120_SLICE_X115Y120_DO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_AMUX = CLBLL_R_X75Y120_SLICE_X115Y120_F7AMUX_O;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B = CLBLL_R_X75Y123_SLICE_X114Y123_BO6;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C = CLBLL_R_X75Y123_SLICE_X114Y123_CO6;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D = CLBLL_R_X75Y123_SLICE_X114Y123_DO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A = CLBLL_R_X75Y123_SLICE_X115Y123_AO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B = CLBLL_R_X75Y123_SLICE_X115Y123_BO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C = CLBLL_R_X75Y123_SLICE_X115Y123_CO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D = CLBLL_R_X75Y123_SLICE_X115Y123_DO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A = CLBLL_R_X75Y124_SLICE_X114Y124_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B = CLBLL_R_X75Y124_SLICE_X114Y124_BO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C = CLBLL_R_X75Y124_SLICE_X114Y124_CO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D = CLBLL_R_X75Y124_SLICE_X114Y124_DO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_BMUX = CLBLL_R_X75Y124_SLICE_X114Y124_F8MUX_O;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A = CLBLL_R_X75Y124_SLICE_X115Y124_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B = CLBLL_R_X75Y124_SLICE_X115Y124_BO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C = CLBLL_R_X75Y124_SLICE_X115Y124_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D = CLBLL_R_X75Y124_SLICE_X115Y124_DO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_AMUX = CLBLL_R_X75Y124_SLICE_X115Y124_F7AMUX_O;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_CMUX = CLBLL_R_X75Y124_SLICE_X115Y124_F7BMUX_O;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_A = CLBLL_R_X75Y125_SLICE_X114Y125_AO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_B = CLBLL_R_X75Y125_SLICE_X114Y125_BO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_C = CLBLL_R_X75Y125_SLICE_X114Y125_CO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_D = CLBLL_R_X75Y125_SLICE_X114Y125_DO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_AMUX = CLBLL_R_X75Y125_SLICE_X114Y125_F7AMUX_O;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_A = CLBLL_R_X75Y125_SLICE_X115Y125_AO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_B = CLBLL_R_X75Y125_SLICE_X115Y125_BO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_C = CLBLL_R_X75Y125_SLICE_X115Y125_CO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_D = CLBLL_R_X75Y125_SLICE_X115Y125_DO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_AMUX = CLBLL_R_X75Y125_SLICE_X115Y125_F7AMUX_O;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_A = CLBLL_R_X75Y126_SLICE_X114Y126_AO6;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_B = CLBLL_R_X75Y126_SLICE_X114Y126_BO6;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_C = CLBLL_R_X75Y126_SLICE_X114Y126_CO6;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_D = CLBLL_R_X75Y126_SLICE_X114Y126_DO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_A = CLBLL_R_X75Y126_SLICE_X115Y126_AO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_B = CLBLL_R_X75Y126_SLICE_X115Y126_BO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_C = CLBLL_R_X75Y126_SLICE_X115Y126_CO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_D = CLBLL_R_X75Y126_SLICE_X115Y126_DO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_AMUX = CLBLL_R_X75Y126_SLICE_X115Y126_F7AMUX_O;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_CMUX = CLBLL_R_X75Y126_SLICE_X115Y126_F7BMUX_O;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A = CLBLL_R_X75Y127_SLICE_X114Y127_AO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B = CLBLL_R_X75Y127_SLICE_X114Y127_BO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C = CLBLL_R_X75Y127_SLICE_X114Y127_CO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D = CLBLL_R_X75Y127_SLICE_X114Y127_DO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_AMUX = CLBLL_R_X75Y127_SLICE_X114Y127_F7AMUX_O;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A = CLBLL_R_X75Y127_SLICE_X115Y127_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B = CLBLL_R_X75Y127_SLICE_X115Y127_BO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C = CLBLL_R_X75Y127_SLICE_X115Y127_CO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D = CLBLL_R_X75Y127_SLICE_X115Y127_DO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_BMUX = CLBLL_R_X75Y127_SLICE_X115Y127_F8MUX_O;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A = CLBLL_R_X75Y128_SLICE_X114Y128_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B = CLBLL_R_X75Y128_SLICE_X114Y128_BO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C = CLBLL_R_X75Y128_SLICE_X114Y128_CO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D = CLBLL_R_X75Y128_SLICE_X114Y128_DO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_BMUX = CLBLL_R_X75Y128_SLICE_X114Y128_F8MUX_O;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A = CLBLL_R_X75Y128_SLICE_X115Y128_AO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B = CLBLL_R_X75Y128_SLICE_X115Y128_BO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D = CLBLL_R_X75Y128_SLICE_X115Y128_DO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_AMUX = CLBLL_R_X75Y128_SLICE_X115Y128_F7AMUX_O;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A = CLBLL_R_X77Y113_SLICE_X119Y113_AO6;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B = CLBLL_R_X77Y113_SLICE_X119Y113_BO6;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C = CLBLL_R_X77Y113_SLICE_X119Y113_CO6;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D = CLBLL_R_X77Y113_SLICE_X119Y113_DO6;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_A = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_B = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_C = CLBLL_R_X77Y114_SLICE_X118Y114_CO6;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_D = CLBLL_R_X77Y114_SLICE_X118Y114_DO6;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_A = CLBLL_R_X77Y114_SLICE_X119Y114_AO6;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_B = CLBLL_R_X77Y114_SLICE_X119Y114_BO6;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_C = CLBLL_R_X77Y114_SLICE_X119Y114_CO6;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_D = CLBLL_R_X77Y114_SLICE_X119Y114_DO6;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_A = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_B = CLBLL_R_X77Y115_SLICE_X118Y115_BO6;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_C = CLBLL_R_X77Y115_SLICE_X118Y115_CO6;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_D = CLBLL_R_X77Y115_SLICE_X118Y115_DO6;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_A = CLBLL_R_X77Y115_SLICE_X119Y115_AO6;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_B = CLBLL_R_X77Y115_SLICE_X119Y115_BO6;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_C = CLBLL_R_X77Y115_SLICE_X119Y115_CO6;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_D = CLBLL_R_X77Y115_SLICE_X119Y115_DO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A = CLBLL_R_X77Y122_SLICE_X119Y122_AO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B = CLBLL_R_X77Y122_SLICE_X119Y122_BO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C = CLBLL_R_X77Y122_SLICE_X119Y122_CO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D = CLBLL_R_X77Y122_SLICE_X119Y122_DO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A = CLBLL_R_X77Y125_SLICE_X118Y125_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B = CLBLL_R_X77Y125_SLICE_X118Y125_BO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C = CLBLL_R_X77Y125_SLICE_X118Y125_CO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D = CLBLL_R_X77Y125_SLICE_X118Y125_DO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_BMUX = CLBLL_R_X77Y125_SLICE_X118Y125_F8MUX_O;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A = CLBLL_R_X77Y125_SLICE_X119Y125_AO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B = CLBLL_R_X77Y125_SLICE_X119Y125_BO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C = CLBLL_R_X77Y125_SLICE_X119Y125_CO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D = CLBLL_R_X77Y125_SLICE_X119Y125_DO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A = CLBLL_R_X77Y129_SLICE_X119Y129_AO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B = CLBLL_R_X77Y129_SLICE_X119Y129_BO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C = CLBLL_R_X77Y129_SLICE_X119Y129_CO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D = CLBLL_R_X77Y129_SLICE_X119Y129_DO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A = CLBLL_R_X77Y130_SLICE_X119Y130_AO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B = CLBLL_R_X77Y130_SLICE_X119Y130_BO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C = CLBLL_R_X77Y130_SLICE_X119Y130_CO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D = CLBLL_R_X77Y130_SLICE_X119Y130_DO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A = CLBLL_R_X77Y131_SLICE_X119Y131_AO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B = CLBLL_R_X77Y131_SLICE_X119Y131_BO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C = CLBLL_R_X77Y131_SLICE_X119Y131_CO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D = CLBLL_R_X77Y131_SLICE_X119Y131_DO6;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_A = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_B = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_C = CLBLL_R_X77Y133_SLICE_X118Y133_CO6;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_D = CLBLL_R_X77Y133_SLICE_X118Y133_DO6;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_A = CLBLL_R_X77Y133_SLICE_X119Y133_AO6;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_B = CLBLL_R_X77Y133_SLICE_X119Y133_BO6;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_C = CLBLL_R_X77Y133_SLICE_X119Y133_CO6;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_D = CLBLL_R_X77Y133_SLICE_X119Y133_DO6;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_A = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_B = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_C = CLBLL_R_X79Y123_SLICE_X122Y123_CO6;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_D = CLBLL_R_X79Y123_SLICE_X122Y123_DO6;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_A = CLBLL_R_X79Y123_SLICE_X123Y123_AO6;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_B = CLBLL_R_X79Y123_SLICE_X123Y123_BO6;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_C = CLBLL_R_X79Y123_SLICE_X123Y123_CO6;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_D = CLBLL_R_X79Y123_SLICE_X123Y123_DO6;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_A = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_B = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_C = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_D = CLBLL_R_X79Y124_SLICE_X122Y124_DO6;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_A = CLBLL_R_X79Y124_SLICE_X123Y124_AO6;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_B = CLBLL_R_X79Y124_SLICE_X123Y124_BO6;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_C = CLBLL_R_X79Y124_SLICE_X123Y124_CO6;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_D = CLBLL_R_X79Y124_SLICE_X123Y124_DO6;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_A = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_B = CLBLL_R_X79Y125_SLICE_X122Y125_BO6;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_C = CLBLL_R_X79Y125_SLICE_X122Y125_CO6;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_D = CLBLL_R_X79Y125_SLICE_X122Y125_DO6;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_A = CLBLL_R_X79Y125_SLICE_X123Y125_AO6;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_B = CLBLL_R_X79Y125_SLICE_X123Y125_BO6;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_C = CLBLL_R_X79Y125_SLICE_X123Y125_CO6;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_D = CLBLL_R_X79Y125_SLICE_X123Y125_DO6;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_A = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_B = CLBLM_L_X44Y118_SLICE_X66Y118_BO6;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_C = CLBLM_L_X44Y118_SLICE_X66Y118_CO6;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_D = CLBLM_L_X44Y118_SLICE_X66Y118_DO6;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_A = CLBLM_L_X44Y118_SLICE_X67Y118_AO6;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_B = CLBLM_L_X44Y118_SLICE_X67Y118_BO6;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_C = CLBLM_L_X44Y118_SLICE_X67Y118_CO6;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_D = CLBLM_L_X44Y118_SLICE_X67Y118_DO6;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_A = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_B = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_C = CLBLM_L_X46Y116_SLICE_X70Y116_CO6;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_D = CLBLM_L_X46Y116_SLICE_X70Y116_DO6;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_A = CLBLM_L_X46Y116_SLICE_X71Y116_AO6;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_B = CLBLM_L_X46Y116_SLICE_X71Y116_BO6;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_C = CLBLM_L_X46Y116_SLICE_X71Y116_CO6;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_D = CLBLM_L_X46Y116_SLICE_X71Y116_DO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_A = CLBLM_L_X56Y116_SLICE_X84Y116_AO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_B = CLBLM_L_X56Y116_SLICE_X84Y116_BO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_C = CLBLM_L_X56Y116_SLICE_X84Y116_CO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_D = CLBLM_L_X56Y116_SLICE_X84Y116_DO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_AMUX = CLBLM_L_X56Y116_SLICE_X84Y116_AO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_CMUX = CLBLM_L_X56Y116_SLICE_X84Y116_CO6;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_A = CLBLM_L_X56Y116_SLICE_X85Y116_AO6;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_B = CLBLM_L_X56Y116_SLICE_X85Y116_BO6;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_C = CLBLM_L_X56Y116_SLICE_X85Y116_CO6;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_D = CLBLM_L_X56Y116_SLICE_X85Y116_DO6;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_A = CLBLM_L_X68Y119_SLICE_X102Y119_AO6;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_B = CLBLM_L_X68Y119_SLICE_X102Y119_BO6;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_C = CLBLM_L_X68Y119_SLICE_X102Y119_CO6;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_D = CLBLM_L_X68Y119_SLICE_X102Y119_DO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_A = CLBLM_L_X68Y119_SLICE_X103Y119_AO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_B = CLBLM_L_X68Y119_SLICE_X103Y119_BO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_C = CLBLM_L_X68Y119_SLICE_X103Y119_CO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_D = CLBLM_L_X68Y119_SLICE_X103Y119_DO6;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_A = CLBLM_L_X70Y117_SLICE_X104Y117_AO6;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_B = CLBLM_L_X70Y117_SLICE_X104Y117_BO6;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_C = CLBLM_L_X70Y117_SLICE_X104Y117_CO6;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_D = CLBLM_L_X70Y117_SLICE_X104Y117_DO6;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_A = CLBLM_L_X70Y117_SLICE_X105Y117_AO6;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_B = CLBLM_L_X70Y117_SLICE_X105Y117_BO6;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_C = CLBLM_L_X70Y117_SLICE_X105Y117_CO6;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_D = CLBLM_L_X70Y117_SLICE_X105Y117_DO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A = CLBLM_L_X70Y119_SLICE_X104Y119_AO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B = CLBLM_L_X70Y119_SLICE_X104Y119_BO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C = CLBLM_L_X70Y119_SLICE_X104Y119_CO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D = CLBLM_L_X70Y119_SLICE_X104Y119_DO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_BMUX = CLBLM_L_X70Y119_SLICE_X104Y119_BO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A = CLBLM_L_X70Y119_SLICE_X105Y119_AO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B = CLBLM_L_X70Y119_SLICE_X105Y119_BO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C = CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D = CLBLM_L_X70Y119_SLICE_X105Y119_DO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_A = CLBLM_L_X70Y121_SLICE_X104Y121_AO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_B = CLBLM_L_X70Y121_SLICE_X104Y121_BO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_C = CLBLM_L_X70Y121_SLICE_X104Y121_CO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_D = CLBLM_L_X70Y121_SLICE_X104Y121_DO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_BMUX = CLBLM_L_X70Y121_SLICE_X104Y121_BO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_CMUX = CLBLM_L_X70Y121_SLICE_X104Y121_CO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_A = CLBLM_L_X70Y121_SLICE_X105Y121_AO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_B = CLBLM_L_X70Y121_SLICE_X105Y121_BO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_C = CLBLM_L_X70Y121_SLICE_X105Y121_CO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_D = CLBLM_L_X70Y121_SLICE_X105Y121_DO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_AMUX = CLBLM_L_X70Y121_SLICE_X105Y121_AO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_BMUX = CLBLM_L_X70Y121_SLICE_X105Y121_BO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_A = CLBLM_L_X70Y122_SLICE_X104Y122_AO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_B = CLBLM_L_X70Y122_SLICE_X104Y122_BO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_C = CLBLM_L_X70Y122_SLICE_X104Y122_CO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_D = CLBLM_L_X70Y122_SLICE_X104Y122_DO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_AMUX = CLBLM_L_X70Y122_SLICE_X104Y122_AO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_CMUX = CLBLM_L_X70Y122_SLICE_X104Y122_CO6;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_A = CLBLM_L_X70Y122_SLICE_X105Y122_AO6;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_B = CLBLM_L_X70Y122_SLICE_X105Y122_BO6;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_C = CLBLM_L_X70Y122_SLICE_X105Y122_CO6;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_D = CLBLM_L_X70Y122_SLICE_X105Y122_DO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A = CLBLM_L_X70Y123_SLICE_X104Y123_AO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B = CLBLM_L_X70Y123_SLICE_X104Y123_BO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C = CLBLM_L_X70Y123_SLICE_X104Y123_CO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D = CLBLM_L_X70Y123_SLICE_X104Y123_DO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A = CLBLM_L_X70Y123_SLICE_X105Y123_AO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B = CLBLM_L_X70Y123_SLICE_X105Y123_BO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C = CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D = CLBLM_L_X70Y123_SLICE_X105Y123_DO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A = CLBLM_L_X70Y124_SLICE_X104Y124_AO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B = CLBLM_L_X70Y124_SLICE_X104Y124_BO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C = CLBLM_L_X70Y124_SLICE_X104Y124_CO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D = CLBLM_L_X70Y124_SLICE_X104Y124_DO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C = CLBLM_L_X70Y124_SLICE_X105Y124_CO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D = CLBLM_L_X70Y124_SLICE_X105Y124_DO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_A = CLBLM_L_X70Y127_SLICE_X104Y127_AO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_B = CLBLM_L_X70Y127_SLICE_X104Y127_BO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_C = CLBLM_L_X70Y127_SLICE_X104Y127_CO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_D = CLBLM_L_X70Y127_SLICE_X104Y127_DO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_AMUX = CLBLM_L_X70Y127_SLICE_X104Y127_AO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_BMUX = CLBLM_L_X70Y127_SLICE_X104Y127_BO6;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_A = CLBLM_L_X70Y127_SLICE_X105Y127_AO6;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_B = CLBLM_L_X70Y127_SLICE_X105Y127_BO6;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_C = CLBLM_L_X70Y127_SLICE_X105Y127_CO6;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_D = CLBLM_L_X70Y127_SLICE_X105Y127_DO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A = CLBLM_L_X70Y128_SLICE_X104Y128_AO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C = CLBLM_L_X70Y128_SLICE_X104Y128_CO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D = CLBLM_L_X70Y128_SLICE_X104Y128_DO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_BMUX = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A = CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B = CLBLM_L_X70Y128_SLICE_X105Y128_BO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C = CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D = CLBLM_L_X70Y128_SLICE_X105Y128_DO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_AMUX = CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A = CLBLM_L_X70Y129_SLICE_X104Y129_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B = CLBLM_L_X70Y129_SLICE_X104Y129_BO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C = CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D = CLBLM_L_X70Y129_SLICE_X104Y129_DO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_AMUX = CLBLM_L_X70Y129_SLICE_X104Y129_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_BMUX = CLBLM_L_X70Y129_SLICE_X104Y129_BO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_CMUX = CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A = CLBLM_L_X70Y129_SLICE_X105Y129_AO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B = CLBLM_L_X70Y129_SLICE_X105Y129_BO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C = CLBLM_L_X70Y129_SLICE_X105Y129_CO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D = CLBLM_L_X70Y129_SLICE_X105Y129_DO6;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_A = CLBLM_L_X72Y114_SLICE_X108Y114_AO6;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_B = CLBLM_L_X72Y114_SLICE_X108Y114_BO6;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_C = CLBLM_L_X72Y114_SLICE_X108Y114_CO6;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_D = CLBLM_L_X72Y114_SLICE_X108Y114_DO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_A = CLBLM_L_X72Y114_SLICE_X109Y114_AO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_B = CLBLM_L_X72Y114_SLICE_X109Y114_BO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_C = CLBLM_L_X72Y114_SLICE_X109Y114_CO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_D = CLBLM_L_X72Y114_SLICE_X109Y114_DO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_AMUX = CLBLM_L_X72Y114_SLICE_X109Y114_F7AMUX_O;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_A = CLBLM_L_X72Y115_SLICE_X108Y115_AO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_B = CLBLM_L_X72Y115_SLICE_X108Y115_BO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_C = CLBLM_L_X72Y115_SLICE_X108Y115_CO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_D = CLBLM_L_X72Y115_SLICE_X108Y115_DO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_BMUX = CLBLM_L_X72Y115_SLICE_X108Y115_F8MUX_O;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_A = CLBLM_L_X72Y115_SLICE_X109Y115_AO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_B = CLBLM_L_X72Y115_SLICE_X109Y115_BO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_C = CLBLM_L_X72Y115_SLICE_X109Y115_CO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_D = CLBLM_L_X72Y115_SLICE_X109Y115_DO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_AMUX = CLBLM_L_X72Y115_SLICE_X109Y115_F7AMUX_O;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_CMUX = CLBLM_L_X72Y115_SLICE_X109Y115_F7BMUX_O;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A = CLBLM_L_X72Y116_SLICE_X108Y116_AO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B = CLBLM_L_X72Y116_SLICE_X108Y116_BO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C = CLBLM_L_X72Y116_SLICE_X108Y116_CO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D = CLBLM_L_X72Y116_SLICE_X108Y116_DO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_AMUX = CLBLM_L_X72Y116_SLICE_X108Y116_F7AMUX_O;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A = CLBLM_L_X72Y116_SLICE_X109Y116_AO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B = CLBLM_L_X72Y116_SLICE_X109Y116_BO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C = CLBLM_L_X72Y116_SLICE_X109Y116_CO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D = CLBLM_L_X72Y116_SLICE_X109Y116_DO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_AMUX = CLBLM_L_X72Y116_SLICE_X109Y116_F7AMUX_O;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_CMUX = CLBLM_L_X72Y116_SLICE_X109Y116_F7BMUX_O;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A = CLBLM_L_X72Y117_SLICE_X108Y117_AO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B = CLBLM_L_X72Y117_SLICE_X108Y117_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C = CLBLM_L_X72Y117_SLICE_X108Y117_CO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D = CLBLM_L_X72Y117_SLICE_X108Y117_DO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_AMUX = CLBLM_L_X72Y117_SLICE_X108Y117_F7AMUX_O;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_CMUX = CLBLM_L_X72Y117_SLICE_X108Y117_F7BMUX_O;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A = CLBLM_L_X72Y117_SLICE_X109Y117_AO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B = CLBLM_L_X72Y117_SLICE_X109Y117_BO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C = CLBLM_L_X72Y117_SLICE_X109Y117_CO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D = CLBLM_L_X72Y117_SLICE_X109Y117_DO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_AMUX = CLBLM_L_X72Y117_SLICE_X109Y117_F7AMUX_O;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A = CLBLM_L_X72Y118_SLICE_X108Y118_AO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B = CLBLM_L_X72Y118_SLICE_X108Y118_BO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C = CLBLM_L_X72Y118_SLICE_X108Y118_CO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D = CLBLM_L_X72Y118_SLICE_X108Y118_DO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_AMUX = CLBLM_L_X72Y118_SLICE_X108Y118_F7AMUX_O;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A = CLBLM_L_X72Y118_SLICE_X109Y118_AO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B = CLBLM_L_X72Y118_SLICE_X109Y118_BO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C = CLBLM_L_X72Y118_SLICE_X109Y118_CO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D = CLBLM_L_X72Y118_SLICE_X109Y118_DO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_AMUX = CLBLM_L_X72Y118_SLICE_X109Y118_F7AMUX_O;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_CMUX = CLBLM_L_X72Y118_SLICE_X109Y118_F7BMUX_O;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A = CLBLM_L_X72Y119_SLICE_X108Y119_AO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B = CLBLM_L_X72Y119_SLICE_X108Y119_BO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C = CLBLM_L_X72Y119_SLICE_X108Y119_CO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D = CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_AMUX = CLBLM_L_X72Y119_SLICE_X108Y119_F7AMUX_O;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A = CLBLM_L_X72Y119_SLICE_X109Y119_AO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B = CLBLM_L_X72Y119_SLICE_X109Y119_BO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C = CLBLM_L_X72Y119_SLICE_X109Y119_CO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D = CLBLM_L_X72Y119_SLICE_X109Y119_DO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_AMUX = CLBLM_L_X72Y119_SLICE_X109Y119_F7AMUX_O;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_CMUX = CLBLM_L_X72Y119_SLICE_X109Y119_F7BMUX_O;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A = CLBLM_L_X72Y120_SLICE_X108Y120_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B = CLBLM_L_X72Y120_SLICE_X108Y120_BO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C = CLBLM_L_X72Y120_SLICE_X108Y120_CO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D = CLBLM_L_X72Y120_SLICE_X108Y120_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_AMUX = CLBLM_L_X72Y120_SLICE_X108Y120_F7AMUX_O;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A = CLBLM_L_X72Y120_SLICE_X109Y120_AO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B = CLBLM_L_X72Y120_SLICE_X109Y120_BO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C = CLBLM_L_X72Y120_SLICE_X109Y120_CO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D = CLBLM_L_X72Y120_SLICE_X109Y120_DO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_BMUX = CLBLM_L_X72Y120_SLICE_X109Y120_F8MUX_O;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A = CLBLM_L_X72Y121_SLICE_X108Y121_AO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B = CLBLM_L_X72Y121_SLICE_X108Y121_BO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C = CLBLM_L_X72Y121_SLICE_X108Y121_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D = CLBLM_L_X72Y121_SLICE_X108Y121_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_BMUX = CLBLM_L_X72Y121_SLICE_X108Y121_F8MUX_O;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A = CLBLM_L_X72Y121_SLICE_X109Y121_AO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B = CLBLM_L_X72Y121_SLICE_X109Y121_BO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C = CLBLM_L_X72Y121_SLICE_X109Y121_CO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D = CLBLM_L_X72Y121_SLICE_X109Y121_DO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_BMUX = CLBLM_L_X72Y121_SLICE_X109Y121_F8MUX_O;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A = CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B = CLBLM_L_X72Y122_SLICE_X108Y122_BO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C = CLBLM_L_X72Y122_SLICE_X108Y122_CO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D = CLBLM_L_X72Y122_SLICE_X108Y122_DO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A = CLBLM_L_X72Y122_SLICE_X109Y122_AO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B = CLBLM_L_X72Y122_SLICE_X109Y122_BO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C = CLBLM_L_X72Y122_SLICE_X109Y122_CO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D = CLBLM_L_X72Y122_SLICE_X109Y122_DO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A = CLBLM_L_X72Y123_SLICE_X108Y123_AO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B = CLBLM_L_X72Y123_SLICE_X108Y123_BO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C = CLBLM_L_X72Y123_SLICE_X108Y123_CO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D = CLBLM_L_X72Y123_SLICE_X108Y123_DO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_AMUX = CLBLM_L_X72Y123_SLICE_X108Y123_F7AMUX_O;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_CMUX = CLBLM_L_X72Y123_SLICE_X108Y123_F7BMUX_O;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A = CLBLM_L_X72Y123_SLICE_X109Y123_AO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B = CLBLM_L_X72Y123_SLICE_X109Y123_BO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C = CLBLM_L_X72Y123_SLICE_X109Y123_CO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D = CLBLM_L_X72Y123_SLICE_X109Y123_DO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_BMUX = CLBLM_L_X72Y123_SLICE_X109Y123_F8MUX_O;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A = CLBLM_L_X72Y124_SLICE_X108Y124_AO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B = CLBLM_L_X72Y124_SLICE_X108Y124_BO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C = CLBLM_L_X72Y124_SLICE_X108Y124_CO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D = CLBLM_L_X72Y124_SLICE_X108Y124_DO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_AMUX = CLBLM_L_X72Y124_SLICE_X108Y124_F7AMUX_O;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A = CLBLM_L_X72Y124_SLICE_X109Y124_AO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B = CLBLM_L_X72Y124_SLICE_X109Y124_BO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C = CLBLM_L_X72Y124_SLICE_X109Y124_CO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D = CLBLM_L_X72Y124_SLICE_X109Y124_DO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_AMUX = CLBLM_L_X72Y124_SLICE_X109Y124_F7AMUX_O;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_CMUX = CLBLM_L_X72Y124_SLICE_X109Y124_F7BMUX_O;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A = CLBLM_L_X72Y125_SLICE_X108Y125_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B = CLBLM_L_X72Y125_SLICE_X108Y125_BO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C = CLBLM_L_X72Y125_SLICE_X108Y125_CO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D = CLBLM_L_X72Y125_SLICE_X108Y125_DO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_AMUX = CLBLM_L_X72Y125_SLICE_X108Y125_F7AMUX_O;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_CMUX = CLBLM_L_X72Y125_SLICE_X108Y125_F7BMUX_O;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A = CLBLM_L_X72Y125_SLICE_X109Y125_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B = CLBLM_L_X72Y125_SLICE_X109Y125_BO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C = CLBLM_L_X72Y125_SLICE_X109Y125_CO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D = CLBLM_L_X72Y125_SLICE_X109Y125_DO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_BMUX = CLBLM_L_X72Y125_SLICE_X109Y125_F8MUX_O;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A = CLBLM_L_X72Y126_SLICE_X108Y126_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B = CLBLM_L_X72Y126_SLICE_X108Y126_BO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C = CLBLM_L_X72Y126_SLICE_X108Y126_CO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D = CLBLM_L_X72Y126_SLICE_X108Y126_DO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_BMUX = CLBLM_L_X72Y126_SLICE_X108Y126_F8MUX_O;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A = CLBLM_L_X72Y126_SLICE_X109Y126_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B = CLBLM_L_X72Y126_SLICE_X109Y126_BO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C = CLBLM_L_X72Y126_SLICE_X109Y126_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D = CLBLM_L_X72Y126_SLICE_X109Y126_DO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_AMUX = CLBLM_L_X72Y126_SLICE_X109Y126_F7AMUX_O;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_CMUX = CLBLM_L_X72Y126_SLICE_X109Y126_F7BMUX_O;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A = CLBLM_L_X72Y127_SLICE_X108Y127_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B = CLBLM_L_X72Y127_SLICE_X108Y127_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C = CLBLM_L_X72Y127_SLICE_X108Y127_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D = CLBLM_L_X72Y127_SLICE_X108Y127_DO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_AMUX = CLBLM_L_X72Y127_SLICE_X108Y127_F7AMUX_O;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_CMUX = CLBLM_L_X72Y127_SLICE_X108Y127_F7BMUX_O;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A = CLBLM_L_X72Y127_SLICE_X109Y127_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B = CLBLM_L_X72Y127_SLICE_X109Y127_BO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C = CLBLM_L_X72Y127_SLICE_X109Y127_CO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D = CLBLM_L_X72Y127_SLICE_X109Y127_DO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_BMUX = CLBLM_L_X72Y127_SLICE_X109Y127_F8MUX_O;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A = CLBLM_L_X72Y128_SLICE_X108Y128_AO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B = CLBLM_L_X72Y128_SLICE_X108Y128_BO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C = CLBLM_L_X72Y128_SLICE_X108Y128_CO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D = CLBLM_L_X72Y128_SLICE_X108Y128_DO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_AMUX = CLBLM_L_X72Y128_SLICE_X108Y128_F7AMUX_O;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A = CLBLM_L_X72Y128_SLICE_X109Y128_AO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B = CLBLM_L_X72Y128_SLICE_X109Y128_BO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C = CLBLM_L_X72Y128_SLICE_X109Y128_CO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D = CLBLM_L_X72Y128_SLICE_X109Y128_DO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_AMUX = CLBLM_L_X72Y128_SLICE_X109Y128_F7AMUX_O;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A = CLBLM_L_X72Y129_SLICE_X108Y129_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B = CLBLM_L_X72Y129_SLICE_X108Y129_BO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C = CLBLM_L_X72Y129_SLICE_X108Y129_CO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D = CLBLM_L_X72Y129_SLICE_X108Y129_DO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_BMUX = CLBLM_L_X72Y129_SLICE_X108Y129_F8MUX_O;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A = CLBLM_L_X72Y129_SLICE_X109Y129_AO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B = CLBLM_L_X72Y129_SLICE_X109Y129_BO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C = CLBLM_L_X72Y129_SLICE_X109Y129_CO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D = CLBLM_L_X72Y129_SLICE_X109Y129_DO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_AMUX = CLBLM_L_X72Y129_SLICE_X109Y129_F7AMUX_O;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_CMUX = CLBLM_L_X72Y129_SLICE_X109Y129_F7BMUX_O;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A = CLBLM_L_X72Y131_SLICE_X108Y131_AO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B = CLBLM_L_X72Y131_SLICE_X108Y131_BO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C = CLBLM_L_X72Y131_SLICE_X108Y131_CO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D = CLBLM_L_X72Y131_SLICE_X108Y131_DO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A = CLBLM_L_X72Y131_SLICE_X109Y131_AO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B = CLBLM_L_X72Y131_SLICE_X109Y131_BO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C = CLBLM_L_X72Y131_SLICE_X109Y131_CO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D = CLBLM_L_X72Y131_SLICE_X109Y131_DO6;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_A = CLBLM_L_X74Y115_SLICE_X112Y115_AO6;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_B = CLBLM_L_X74Y115_SLICE_X112Y115_BO6;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_C = CLBLM_L_X74Y115_SLICE_X112Y115_CO6;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_D = CLBLM_L_X74Y115_SLICE_X112Y115_DO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_A = CLBLM_L_X74Y115_SLICE_X113Y115_AO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_B = CLBLM_L_X74Y115_SLICE_X113Y115_BO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_C = CLBLM_L_X74Y115_SLICE_X113Y115_CO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_D = CLBLM_L_X74Y115_SLICE_X113Y115_DO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_BMUX = CLBLM_L_X74Y115_SLICE_X113Y115_F8MUX_O;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_A = CLBLM_L_X74Y116_SLICE_X112Y116_AO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_B = CLBLM_L_X74Y116_SLICE_X112Y116_BO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_C = CLBLM_L_X74Y116_SLICE_X112Y116_CO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_D = CLBLM_L_X74Y116_SLICE_X112Y116_DO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_BMUX = CLBLM_L_X74Y116_SLICE_X112Y116_F8MUX_O;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_A = CLBLM_L_X74Y116_SLICE_X113Y116_AO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_B = CLBLM_L_X74Y116_SLICE_X113Y116_BO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_C = CLBLM_L_X74Y116_SLICE_X113Y116_CO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_D = CLBLM_L_X74Y116_SLICE_X113Y116_DO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_AMUX = CLBLM_L_X74Y116_SLICE_X113Y116_F7AMUX_O;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A = CLBLM_L_X74Y117_SLICE_X112Y117_AO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B = CLBLM_L_X74Y117_SLICE_X112Y117_BO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C = CLBLM_L_X74Y117_SLICE_X112Y117_CO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D = CLBLM_L_X74Y117_SLICE_X112Y117_DO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_BMUX = CLBLM_L_X74Y117_SLICE_X112Y117_F8MUX_O;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A = CLBLM_L_X74Y117_SLICE_X113Y117_AO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B = CLBLM_L_X74Y117_SLICE_X113Y117_BO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C = CLBLM_L_X74Y117_SLICE_X113Y117_CO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D = CLBLM_L_X74Y117_SLICE_X113Y117_DO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_AMUX = CLBLM_L_X74Y117_SLICE_X113Y117_F7AMUX_O;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A = CLBLM_L_X74Y118_SLICE_X112Y118_AO6;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B = CLBLM_L_X74Y118_SLICE_X112Y118_BO6;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C = CLBLM_L_X74Y118_SLICE_X112Y118_CO6;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D = CLBLM_L_X74Y118_SLICE_X112Y118_DO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A = CLBLM_L_X74Y118_SLICE_X113Y118_AO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B = CLBLM_L_X74Y118_SLICE_X113Y118_BO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C = CLBLM_L_X74Y118_SLICE_X113Y118_CO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D = CLBLM_L_X74Y118_SLICE_X113Y118_DO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_AMUX = CLBLM_L_X74Y118_SLICE_X113Y118_F7AMUX_O;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A = CLBLM_L_X74Y119_SLICE_X112Y119_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B = CLBLM_L_X74Y119_SLICE_X112Y119_BO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C = CLBLM_L_X74Y119_SLICE_X112Y119_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D = CLBLM_L_X74Y119_SLICE_X112Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_BMUX = CLBLM_L_X74Y119_SLICE_X112Y119_F8MUX_O;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A = CLBLM_L_X74Y119_SLICE_X113Y119_AO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B = CLBLM_L_X74Y119_SLICE_X113Y119_BO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C = CLBLM_L_X74Y119_SLICE_X113Y119_CO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D = CLBLM_L_X74Y119_SLICE_X113Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_AMUX = CLBLM_L_X74Y119_SLICE_X113Y119_F7AMUX_O;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_CMUX = CLBLM_L_X74Y119_SLICE_X113Y119_F7BMUX_O;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A = CLBLM_L_X74Y120_SLICE_X112Y120_AO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B = CLBLM_L_X74Y120_SLICE_X112Y120_BO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C = CLBLM_L_X74Y120_SLICE_X112Y120_CO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D = CLBLM_L_X74Y120_SLICE_X112Y120_DO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_BMUX = CLBLM_L_X74Y120_SLICE_X112Y120_F8MUX_O;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A = CLBLM_L_X74Y120_SLICE_X113Y120_AO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B = CLBLM_L_X74Y120_SLICE_X113Y120_BO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C = CLBLM_L_X74Y120_SLICE_X113Y120_CO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D = CLBLM_L_X74Y120_SLICE_X113Y120_DO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_AMUX = CLBLM_L_X74Y120_SLICE_X113Y120_AO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A = CLBLM_L_X74Y121_SLICE_X112Y121_AO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B = CLBLM_L_X74Y121_SLICE_X112Y121_BO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C = CLBLM_L_X74Y121_SLICE_X112Y121_CO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D = CLBLM_L_X74Y121_SLICE_X112Y121_DO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_BMUX = CLBLM_L_X74Y121_SLICE_X112Y121_F8MUX_O;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A = CLBLM_L_X74Y121_SLICE_X113Y121_AO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B = CLBLM_L_X74Y121_SLICE_X113Y121_BO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C = CLBLM_L_X74Y121_SLICE_X113Y121_CO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D = CLBLM_L_X74Y121_SLICE_X113Y121_DO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_BMUX = CLBLM_L_X74Y121_SLICE_X113Y121_F8MUX_O;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A = CLBLM_L_X74Y123_SLICE_X112Y123_AO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B = CLBLM_L_X74Y123_SLICE_X112Y123_BO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C = CLBLM_L_X74Y123_SLICE_X112Y123_CO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D = CLBLM_L_X74Y123_SLICE_X112Y123_DO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_AMUX = CLBLM_L_X74Y123_SLICE_X112Y123_F7AMUX_O;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A = CLBLM_L_X74Y123_SLICE_X113Y123_AO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B = CLBLM_L_X74Y123_SLICE_X113Y123_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C = CLBLM_L_X74Y123_SLICE_X113Y123_CO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D = CLBLM_L_X74Y123_SLICE_X113Y123_DO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_BMUX = CLBLM_L_X74Y123_SLICE_X113Y123_F8MUX_O;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_A = CLBLM_L_X74Y124_SLICE_X112Y124_AO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_B = CLBLM_L_X74Y124_SLICE_X112Y124_BO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_C = CLBLM_L_X74Y124_SLICE_X112Y124_CO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_D = CLBLM_L_X74Y124_SLICE_X112Y124_DO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_BMUX = CLBLM_L_X74Y124_SLICE_X112Y124_F8MUX_O;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_A = CLBLM_L_X74Y124_SLICE_X113Y124_AO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_B = CLBLM_L_X74Y124_SLICE_X113Y124_BO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_C = CLBLM_L_X74Y124_SLICE_X113Y124_CO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_D = CLBLM_L_X74Y124_SLICE_X113Y124_DO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_AMUX = CLBLM_L_X74Y124_SLICE_X113Y124_F7AMUX_O;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_CMUX = CLBLM_L_X74Y124_SLICE_X113Y124_F7BMUX_O;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A = CLBLM_L_X74Y125_SLICE_X112Y125_AO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B = CLBLM_L_X74Y125_SLICE_X112Y125_BO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C = CLBLM_L_X74Y125_SLICE_X112Y125_CO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D = CLBLM_L_X74Y125_SLICE_X112Y125_DO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_AMUX = CLBLM_L_X74Y125_SLICE_X112Y125_F7AMUX_O;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A = CLBLM_L_X74Y125_SLICE_X113Y125_AO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B = CLBLM_L_X74Y125_SLICE_X113Y125_BO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C = CLBLM_L_X74Y125_SLICE_X113Y125_CO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D = CLBLM_L_X74Y125_SLICE_X113Y125_DO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_AMUX = CLBLM_L_X74Y125_SLICE_X113Y125_F7AMUX_O;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_CMUX = CLBLM_L_X74Y125_SLICE_X113Y125_F7BMUX_O;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A = CLBLM_L_X74Y126_SLICE_X112Y126_AO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B = CLBLM_L_X74Y126_SLICE_X112Y126_BO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C = CLBLM_L_X74Y126_SLICE_X112Y126_CO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D = CLBLM_L_X74Y126_SLICE_X112Y126_DO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_BMUX = CLBLM_L_X74Y126_SLICE_X112Y126_F8MUX_O;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A = CLBLM_L_X74Y126_SLICE_X113Y126_AO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B = CLBLM_L_X74Y126_SLICE_X113Y126_BO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C = CLBLM_L_X74Y126_SLICE_X113Y126_CO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D = CLBLM_L_X74Y126_SLICE_X113Y126_DO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A = CLBLM_L_X74Y127_SLICE_X112Y127_AO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B = CLBLM_L_X74Y127_SLICE_X112Y127_BO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C = CLBLM_L_X74Y127_SLICE_X112Y127_CO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D = CLBLM_L_X74Y127_SLICE_X112Y127_DO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_AMUX = CLBLM_L_X74Y127_SLICE_X112Y127_F7AMUX_O;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_CMUX = CLBLM_L_X74Y127_SLICE_X112Y127_F7BMUX_O;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A = CLBLM_L_X74Y127_SLICE_X113Y127_AO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B = CLBLM_L_X74Y127_SLICE_X113Y127_BO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C = CLBLM_L_X74Y127_SLICE_X113Y127_CO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D = CLBLM_L_X74Y127_SLICE_X113Y127_DO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_AMUX = CLBLM_L_X74Y127_SLICE_X113Y127_F7AMUX_O;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A = CLBLM_L_X74Y128_SLICE_X112Y128_AO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B = CLBLM_L_X74Y128_SLICE_X112Y128_BO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C = CLBLM_L_X74Y128_SLICE_X112Y128_CO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D = CLBLM_L_X74Y128_SLICE_X112Y128_DO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_AMUX = CLBLM_L_X74Y128_SLICE_X112Y128_F7AMUX_O;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A = CLBLM_L_X74Y128_SLICE_X113Y128_AO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B = CLBLM_L_X74Y128_SLICE_X113Y128_BO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C = CLBLM_L_X74Y128_SLICE_X113Y128_CO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D = CLBLM_L_X74Y128_SLICE_X113Y128_DO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_BMUX = CLBLM_L_X74Y128_SLICE_X113Y128_F8MUX_O;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A = CLBLM_L_X74Y129_SLICE_X112Y129_AO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B = CLBLM_L_X74Y129_SLICE_X112Y129_BO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C = CLBLM_L_X74Y129_SLICE_X112Y129_CO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D = CLBLM_L_X74Y129_SLICE_X112Y129_DO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_AMUX = CLBLM_L_X74Y129_SLICE_X112Y129_F7AMUX_O;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A = CLBLM_L_X74Y129_SLICE_X113Y129_AO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B = CLBLM_L_X74Y129_SLICE_X113Y129_BO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C = CLBLM_L_X74Y129_SLICE_X113Y129_CO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D = CLBLM_L_X74Y129_SLICE_X113Y129_DO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_A = CLBLM_L_X76Y120_SLICE_X116Y120_AO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_B = CLBLM_L_X76Y120_SLICE_X116Y120_BO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_C = CLBLM_L_X76Y120_SLICE_X116Y120_CO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_D = CLBLM_L_X76Y120_SLICE_X116Y120_DO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_BMUX = CLBLM_L_X76Y120_SLICE_X116Y120_F8MUX_O;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_A = CLBLM_L_X76Y120_SLICE_X117Y120_AO6;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_B = CLBLM_L_X76Y120_SLICE_X117Y120_BO6;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_C = CLBLM_L_X76Y120_SLICE_X117Y120_CO6;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_D = CLBLM_L_X76Y120_SLICE_X117Y120_DO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A = CLBLM_L_X76Y124_SLICE_X116Y124_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B = CLBLM_L_X76Y124_SLICE_X116Y124_BO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C = CLBLM_L_X76Y124_SLICE_X116Y124_CO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D = CLBLM_L_X76Y124_SLICE_X116Y124_DO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_AMUX = CLBLM_L_X76Y124_SLICE_X116Y124_F7AMUX_O;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_CMUX = CLBLM_L_X76Y124_SLICE_X116Y124_F7BMUX_O;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A = CLBLM_L_X76Y124_SLICE_X117Y124_AO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B = CLBLM_L_X76Y124_SLICE_X117Y124_BO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C = CLBLM_L_X76Y124_SLICE_X117Y124_CO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D = CLBLM_L_X76Y124_SLICE_X117Y124_DO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A = CLBLM_L_X76Y125_SLICE_X116Y125_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B = CLBLM_L_X76Y125_SLICE_X116Y125_BO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C = CLBLM_L_X76Y125_SLICE_X116Y125_CO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D = CLBLM_L_X76Y125_SLICE_X116Y125_DO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_BMUX = CLBLM_L_X76Y125_SLICE_X116Y125_F8MUX_O;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A = CLBLM_L_X76Y125_SLICE_X117Y125_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B = CLBLM_L_X76Y125_SLICE_X117Y125_BO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C = CLBLM_L_X76Y125_SLICE_X117Y125_CO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D = CLBLM_L_X76Y125_SLICE_X117Y125_DO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_BMUX = CLBLM_L_X76Y125_SLICE_X117Y125_F8MUX_O;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A = CLBLM_L_X76Y127_SLICE_X116Y127_AO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B = CLBLM_L_X76Y127_SLICE_X116Y127_BO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D = CLBLM_L_X76Y127_SLICE_X116Y127_DO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_AMUX = CLBLM_L_X76Y127_SLICE_X116Y127_F7AMUX_O;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A = CLBLM_L_X76Y127_SLICE_X117Y127_AO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B = CLBLM_L_X76Y127_SLICE_X117Y127_BO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C = CLBLM_L_X76Y127_SLICE_X117Y127_CO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D = CLBLM_L_X76Y127_SLICE_X117Y127_DO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A = CLBLM_L_X76Y128_SLICE_X116Y128_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B = CLBLM_L_X76Y128_SLICE_X116Y128_BO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C = CLBLM_L_X76Y128_SLICE_X116Y128_CO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D = CLBLM_L_X76Y128_SLICE_X116Y128_DO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_BMUX = CLBLM_L_X76Y128_SLICE_X116Y128_F8MUX_O;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A = CLBLM_L_X76Y128_SLICE_X117Y128_AO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B = CLBLM_L_X76Y128_SLICE_X117Y128_BO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C = CLBLM_L_X76Y128_SLICE_X117Y128_CO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D = CLBLM_L_X76Y128_SLICE_X117Y128_DO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_A = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_B = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_C = CLBLM_L_X76Y131_SLICE_X116Y131_CO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_D = CLBLM_L_X76Y131_SLICE_X116Y131_DO6;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_A = CLBLM_L_X76Y131_SLICE_X117Y131_AO6;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_B = CLBLM_L_X76Y131_SLICE_X117Y131_BO6;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_C = CLBLM_L_X76Y131_SLICE_X117Y131_CO6;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_D = CLBLM_L_X76Y131_SLICE_X117Y131_DO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A = CLBLM_L_X76Y133_SLICE_X116Y133_AO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B = CLBLM_L_X76Y133_SLICE_X116Y133_BO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C = CLBLM_L_X76Y133_SLICE_X116Y133_CO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D = CLBLM_L_X76Y133_SLICE_X116Y133_DO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B = CLBLM_L_X76Y133_SLICE_X117Y133_BO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C = CLBLM_L_X76Y133_SLICE_X117Y133_CO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D = CLBLM_L_X76Y133_SLICE_X117Y133_DO6;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_A = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_B = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_C = CLBLM_L_X78Y117_SLICE_X120Y117_CO6;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_D = CLBLM_L_X78Y117_SLICE_X120Y117_DO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_A = CLBLM_L_X78Y117_SLICE_X121Y117_AO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_B = CLBLM_L_X78Y117_SLICE_X121Y117_BO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_C = CLBLM_L_X78Y117_SLICE_X121Y117_CO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_D = CLBLM_L_X78Y117_SLICE_X121Y117_DO6;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D = CLBLM_L_X78Y119_SLICE_X120Y119_DO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A = CLBLM_L_X78Y119_SLICE_X121Y119_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B = CLBLM_L_X78Y119_SLICE_X121Y119_BO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C = CLBLM_L_X78Y119_SLICE_X121Y119_CO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D = CLBLM_L_X78Y119_SLICE_X121Y119_DO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D = CLBLM_L_X78Y120_SLICE_X120Y120_DO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A = CLBLM_L_X78Y120_SLICE_X121Y120_AO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B = CLBLM_L_X78Y120_SLICE_X121Y120_BO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C = CLBLM_L_X78Y120_SLICE_X121Y120_CO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D = CLBLM_L_X78Y120_SLICE_X121Y120_DO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B = CLBLM_L_X78Y121_SLICE_X120Y121_BO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C = CLBLM_L_X78Y121_SLICE_X120Y121_CO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D = CLBLM_L_X78Y121_SLICE_X120Y121_DO6;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A = CLBLM_L_X78Y121_SLICE_X121Y121_AO6;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B = CLBLM_L_X78Y121_SLICE_X121Y121_BO6;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C = CLBLM_L_X78Y121_SLICE_X121Y121_CO6;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D = CLBLM_L_X78Y121_SLICE_X121Y121_DO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C = CLBLM_L_X78Y122_SLICE_X120Y122_CO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D = CLBLM_L_X78Y122_SLICE_X120Y122_DO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A = CLBLM_L_X78Y122_SLICE_X121Y122_AO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B = CLBLM_L_X78Y122_SLICE_X121Y122_BO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C = CLBLM_L_X78Y122_SLICE_X121Y122_CO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D = CLBLM_L_X78Y122_SLICE_X121Y122_DO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A = CLBLM_L_X78Y123_SLICE_X121Y123_AO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B = CLBLM_L_X78Y123_SLICE_X121Y123_BO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C = CLBLM_L_X78Y123_SLICE_X121Y123_CO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D = CLBLM_L_X78Y123_SLICE_X121Y123_DO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C = CLBLM_L_X78Y124_SLICE_X120Y124_CO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D = CLBLM_L_X78Y124_SLICE_X120Y124_DO6;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A = CLBLM_L_X78Y124_SLICE_X121Y124_AO6;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B = CLBLM_L_X78Y124_SLICE_X121Y124_BO6;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C = CLBLM_L_X78Y124_SLICE_X121Y124_CO6;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D = CLBLM_L_X78Y124_SLICE_X121Y124_DO6;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_A = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_B = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_C = CLBLM_L_X78Y126_SLICE_X120Y126_CO6;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_D = CLBLM_L_X78Y126_SLICE_X120Y126_DO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_A = CLBLM_L_X78Y126_SLICE_X121Y126_AO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_B = CLBLM_L_X78Y126_SLICE_X121Y126_BO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_C = CLBLM_L_X78Y126_SLICE_X121Y126_CO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_D = CLBLM_L_X78Y126_SLICE_X121Y126_DO6;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B = CLBLM_L_X78Y129_SLICE_X120Y129_BO6;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C = CLBLM_L_X78Y129_SLICE_X120Y129_CO6;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D = CLBLM_L_X78Y129_SLICE_X120Y129_DO6;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A = CLBLM_L_X78Y129_SLICE_X121Y129_AO6;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B = CLBLM_L_X78Y129_SLICE_X121Y129_BO6;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C = CLBLM_L_X78Y129_SLICE_X121Y129_CO6;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D = CLBLM_L_X78Y129_SLICE_X121Y129_DO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B = CLBLM_L_X98Y131_SLICE_X154Y131_BO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C = CLBLM_L_X98Y131_SLICE_X154Y131_CO6;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D = CLBLM_L_X98Y131_SLICE_X154Y131_DO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A = CLBLM_L_X98Y131_SLICE_X155Y131_AO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B = CLBLM_L_X98Y131_SLICE_X155Y131_BO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C = CLBLM_L_X98Y131_SLICE_X155Y131_CO6;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D = CLBLM_L_X98Y131_SLICE_X155Y131_DO6;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B = CLBLM_L_X98Y132_SLICE_X154Y132_BO6;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C = CLBLM_L_X98Y132_SLICE_X154Y132_CO6;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D = CLBLM_L_X98Y132_SLICE_X154Y132_DO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A = CLBLM_L_X98Y132_SLICE_X155Y132_AO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B = CLBLM_L_X98Y132_SLICE_X155Y132_BO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C = CLBLM_L_X98Y132_SLICE_X155Y132_CO6;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D = CLBLM_L_X98Y132_SLICE_X155Y132_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_AMUX = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_AMUX = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_A = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_B = CLBLM_R_X49Y116_SLICE_X74Y116_BO6;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_C = CLBLM_R_X49Y116_SLICE_X74Y116_CO6;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_D = CLBLM_R_X49Y116_SLICE_X74Y116_DO6;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_A = CLBLM_R_X49Y116_SLICE_X75Y116_AO6;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_B = CLBLM_R_X49Y116_SLICE_X75Y116_BO6;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_C = CLBLM_R_X49Y116_SLICE_X75Y116_CO6;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_D = CLBLM_R_X49Y116_SLICE_X75Y116_DO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_A = CLBLM_R_X59Y117_SLICE_X88Y117_AO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_B = CLBLM_R_X59Y117_SLICE_X88Y117_BO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_C = CLBLM_R_X59Y117_SLICE_X88Y117_CO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_D = CLBLM_R_X59Y117_SLICE_X88Y117_DO6;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_A = CLBLM_R_X59Y117_SLICE_X89Y117_AO6;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_B = CLBLM_R_X59Y117_SLICE_X89Y117_BO6;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_C = CLBLM_R_X59Y117_SLICE_X89Y117_CO6;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_D = CLBLM_R_X59Y117_SLICE_X89Y117_DO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_A = CLBLM_R_X59Y118_SLICE_X88Y118_AO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_B = CLBLM_R_X59Y118_SLICE_X88Y118_BO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_C = CLBLM_R_X59Y118_SLICE_X88Y118_CO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_D = CLBLM_R_X59Y118_SLICE_X88Y118_DO6;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_A = CLBLM_R_X59Y118_SLICE_X89Y118_AO6;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_B = CLBLM_R_X59Y118_SLICE_X89Y118_BO6;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_C = CLBLM_R_X59Y118_SLICE_X89Y118_CO6;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_D = CLBLM_R_X59Y118_SLICE_X89Y118_DO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_O = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_O = LIOB33_X0Y83_IOB_X0Y84_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_O = LIOB33_X0Y83_IOB_X0Y83_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_O = LIOB33_X0Y85_IOB_X0Y85_I;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_OQ = CLBLM_L_X70Y119_SLICE_X104Y119_AO6;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_TQ = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_OQ = CLBLL_R_X71Y128_SLICE_X106Y128_AO6;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_TQ = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_OQ = CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_TQ = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_OQ = CLBLL_R_X71Y131_SLICE_X107Y131_BO6;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_TQ = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_OQ = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_TQ = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_OQ = CLBLM_L_X70Y124_SLICE_X104Y124_AO6;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_TQ = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_OQ = CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_TQ = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_OQ = CLBLL_R_X71Y131_SLICE_X106Y131_AO6;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_TQ = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_OQ = CLBLM_L_X70Y124_SLICE_X104Y124_CO6;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLM_R_X59Y117_SLICE_X88Y117_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLM_L_X56Y116_SLICE_X84Y116_AO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_L_X70Y123_SLICE_X105Y123_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLM_L_X70Y123_SLICE_X104Y123_BO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_L_X72Y131_SLICE_X108Y131_AO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X70Y121_SLICE_X105Y121_AO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_L_X70Y122_SLICE_X104Y122_CO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_L_X70Y119_SLICE_X105Y119_AO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_L_X70Y121_SLICE_X105Y121_CO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_L_X70Y127_SLICE_X104Y127_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X70Y121_SLICE_X104Y121_DO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_L_X70Y123_SLICE_X105Y123_DO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_L_X70Y127_SLICE_X104Y127_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_L_X70Y127_SLICE_X104Y127_DO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_O = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_O = LIOB33_X0Y151_IOB_X0Y151_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_O = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_O = LIOB33_X0Y153_IOB_X0Y153_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_O = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_O = LIOB33_X0Y155_IOB_X0Y155_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_O = LIOB33_X0Y159_IOB_X0Y160_I;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_O = LIOB33_X0Y159_IOB_X0Y159_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_O = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_O = LIOB33_X0Y161_IOB_X0Y161_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_O = LIOB33_X0Y165_IOB_X0Y166_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_O = LIOB33_X0Y165_IOB_X0Y165_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_O = LIOB33_X0Y167_IOB_X0Y168_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y167_O = LIOB33_X0Y167_IOB_X0Y167_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_O = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_O = LIOB33_X0Y171_IOB_X0Y171_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_O = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_O = LIOB33_X0Y173_IOB_X0Y173_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_O = LIOB33_X0Y175_IOB_X0Y176_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_O = LIOB33_X0Y175_IOB_X0Y175_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_O = LIOB33_X0Y177_IOB_X0Y178_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_O = LIOB33_X0Y177_IOB_X0Y177_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_O = LIOB33_X0Y179_IOB_X0Y180_I;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_O = LIOB33_X0Y179_IOB_X0Y179_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_O = LIOB33_X0Y183_IOB_X0Y184_I;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_O = LIOB33_X0Y183_IOB_X0Y183_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_O = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_O = LIOB33_X0Y185_IOB_X0Y185_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_O = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_O = LIOB33_X0Y189_IOB_X0Y189_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_O = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_O = LIOB33_X0Y191_IOB_X0Y191_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_O = LIOB33_X0Y195_IOB_X0Y196_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_O = LIOB33_X0Y195_IOB_X0Y195_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y198_O = LIOB33_X0Y197_IOB_X0Y198_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_O = LIOB33_X0Y197_IOB_X0Y197_I;
  assign LIOI3_X0Y201_ILOGIC_X0Y202_O = LIOB33_X0Y201_IOB_X0Y202_I;
  assign LIOI3_X0Y201_ILOGIC_X0Y201_O = LIOB33_X0Y201_IOB_X0Y201_I;
  assign LIOI3_X0Y203_ILOGIC_X0Y203_O = LIOB33_X0Y203_IOB_X0Y203_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_OQ = CLBLL_R_X71Y131_SLICE_X106Y131_CO6;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLM_R_X59Y118_SLICE_X88Y118_AO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_O = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign LIOI3_SING_X0Y199_ILOGIC_X0Y199_O = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign LIOI3_SING_X0Y200_ILOGIC_X0Y200_O = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_O = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_O = LIOB33_X0Y81_IOB_X0Y81_I;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_OQ = CLBLM_L_X70Y129_SLICE_X104Y129_AO6;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_OQ = CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLM_L_X70Y121_SLICE_X104Y121_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLM_L_X56Y116_SLICE_X84Y116_CO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_L_X70Y121_SLICE_X104Y121_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_O = LIOB33_X0Y157_IOB_X0Y158_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_O = LIOB33_X0Y157_IOB_X0Y157_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_O = LIOB33_X0Y169_IOB_X0Y170_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_O = LIOB33_X0Y169_IOB_X0Y169_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_O = LIOB33_X0Y181_IOB_X0Y182_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_O = LIOB33_X0Y181_IOB_X0Y181_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_O = LIOB33_X0Y193_IOB_X0Y194_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_O = LIOB33_X0Y193_IOB_X0Y193_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_OQ = CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_OQ = CLBLL_R_X71Y119_SLICE_X106Y119_AO6;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_L_X70Y122_SLICE_X104Y122_AO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_O = LIOB33_X0Y163_IOB_X0Y164_I;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_O = LIOB33_X0Y163_IOB_X0Y163_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_O = LIOB33_X0Y187_IOB_X0Y188_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_O = LIOB33_X0Y187_IOB_X0Y187_I;
  assign RIOI3_X105Y51_ILOGIC_X1Y52_O = RIOB33_X105Y51_IOB_X1Y52_I;
  assign RIOI3_X105Y51_ILOGIC_X1Y51_O = RIOB33_X105Y51_IOB_X1Y51_I;
  assign RIOI3_X105Y53_ILOGIC_X1Y54_O = RIOB33_X105Y53_IOB_X1Y54_I;
  assign RIOI3_X105Y53_ILOGIC_X1Y53_O = RIOB33_X105Y53_IOB_X1Y53_I;
  assign RIOI3_X105Y55_ILOGIC_X1Y56_O = RIOB33_X105Y55_IOB_X1Y56_I;
  assign RIOI3_X105Y55_ILOGIC_X1Y55_O = RIOB33_X105Y55_IOB_X1Y55_I;
  assign RIOI3_X105Y59_ILOGIC_X1Y60_O = RIOB33_X105Y59_IOB_X1Y60_I;
  assign RIOI3_X105Y59_ILOGIC_X1Y59_O = RIOB33_X105Y59_IOB_X1Y59_I;
  assign RIOI3_X105Y61_ILOGIC_X1Y62_O = RIOB33_X105Y61_IOB_X1Y62_I;
  assign RIOI3_X105Y61_ILOGIC_X1Y61_O = RIOB33_X105Y61_IOB_X1Y61_I;
  assign RIOI3_X105Y65_ILOGIC_X1Y66_O = RIOB33_X105Y65_IOB_X1Y66_I;
  assign RIOI3_X105Y65_ILOGIC_X1Y65_O = RIOB33_X105Y65_IOB_X1Y65_I;
  assign RIOI3_X105Y67_ILOGIC_X1Y68_O = RIOB33_X105Y67_IOB_X1Y68_I;
  assign RIOI3_X105Y67_ILOGIC_X1Y67_O = RIOB33_X105Y67_IOB_X1Y67_I;
  assign RIOI3_X105Y71_ILOGIC_X1Y72_O = RIOB33_X105Y71_IOB_X1Y72_I;
  assign RIOI3_X105Y71_ILOGIC_X1Y71_O = RIOB33_X105Y71_IOB_X1Y71_I;
  assign RIOI3_X105Y73_ILOGIC_X1Y74_O = RIOB33_X105Y73_IOB_X1Y74_I;
  assign RIOI3_X105Y73_ILOGIC_X1Y73_O = RIOB33_X105Y73_IOB_X1Y73_I;
  assign RIOI3_X105Y75_ILOGIC_X1Y76_O = RIOB33_X105Y75_IOB_X1Y76_I;
  assign RIOI3_X105Y75_ILOGIC_X1Y75_O = RIOB33_X105Y75_IOB_X1Y75_I;
  assign RIOI3_X105Y77_ILOGIC_X1Y78_O = RIOB33_X105Y77_IOB_X1Y78_I;
  assign RIOI3_X105Y77_ILOGIC_X1Y77_O = RIOB33_X105Y77_IOB_X1Y77_I;
  assign RIOI3_X105Y79_ILOGIC_X1Y80_O = RIOB33_X105Y79_IOB_X1Y80_I;
  assign RIOI3_X105Y79_ILOGIC_X1Y79_O = RIOB33_X105Y79_IOB_X1Y79_I;
  assign RIOI3_X105Y83_ILOGIC_X1Y84_O = RIOB33_X105Y83_IOB_X1Y84_I;
  assign RIOI3_X105Y83_ILOGIC_X1Y83_O = RIOB33_X105Y83_IOB_X1Y83_I;
  assign RIOI3_X105Y85_ILOGIC_X1Y86_O = RIOB33_X105Y85_IOB_X1Y86_I;
  assign RIOI3_X105Y85_ILOGIC_X1Y85_O = RIOB33_X105Y85_IOB_X1Y85_I;
  assign RIOI3_X105Y89_ILOGIC_X1Y90_O = RIOB33_X105Y89_IOB_X1Y90_I;
  assign RIOI3_X105Y89_ILOGIC_X1Y89_O = RIOB33_X105Y89_IOB_X1Y89_I;
  assign RIOI3_X105Y91_ILOGIC_X1Y92_O = RIOB33_X105Y91_IOB_X1Y92_I;
  assign RIOI3_X105Y91_ILOGIC_X1Y91_O = RIOB33_X105Y91_IOB_X1Y91_I;
  assign RIOI3_X105Y95_ILOGIC_X1Y96_O = RIOB33_X105Y95_IOB_X1Y96_I;
  assign RIOI3_X105Y95_ILOGIC_X1Y95_O = RIOB33_X105Y95_IOB_X1Y95_I;
  assign RIOI3_X105Y97_ILOGIC_X1Y98_O = RIOB33_X105Y97_IOB_X1Y98_I;
  assign RIOI3_X105Y97_ILOGIC_X1Y97_O = RIOB33_X105Y97_IOB_X1Y97_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y152_O = RIOB33_X105Y151_IOB_X1Y152_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y151_O = RIOB33_X105Y151_IOB_X1Y151_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y154_O = RIOB33_X105Y153_IOB_X1Y154_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y153_O = RIOB33_X105Y153_IOB_X1Y153_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y156_O = RIOB33_X105Y155_IOB_X1Y156_I;
  assign RIOI3_X105Y155_ILOGIC_X1Y155_O = RIOB33_X105Y155_IOB_X1Y155_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y160_O = RIOB33_X105Y159_IOB_X1Y160_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y159_O = RIOB33_X105Y159_IOB_X1Y159_I;
  assign RIOI3_X105Y161_ILOGIC_X1Y162_O = RIOB33_X105Y161_IOB_X1Y162_I;
  assign RIOI3_X105Y161_ILOGIC_X1Y161_O = RIOB33_X105Y161_IOB_X1Y161_I;
  assign RIOI3_X105Y165_ILOGIC_X1Y166_O = RIOB33_X105Y165_IOB_X1Y166_I;
  assign RIOI3_X105Y165_ILOGIC_X1Y165_O = RIOB33_X105Y165_IOB_X1Y165_I;
  assign RIOI3_X105Y167_ILOGIC_X1Y168_O = RIOB33_X105Y167_IOB_X1Y168_I;
  assign RIOI3_X105Y167_ILOGIC_X1Y167_O = RIOB33_X105Y167_IOB_X1Y167_I;
  assign RIOI3_X105Y171_ILOGIC_X1Y172_O = RIOB33_X105Y171_IOB_X1Y172_I;
  assign RIOI3_X105Y171_ILOGIC_X1Y171_O = RIOB33_X105Y171_IOB_X1Y171_I;
  assign RIOI3_X105Y173_ILOGIC_X1Y174_O = RIOB33_X105Y173_IOB_X1Y174_I;
  assign RIOI3_X105Y173_ILOGIC_X1Y173_O = RIOB33_X105Y173_IOB_X1Y173_I;
  assign RIOI3_X105Y175_ILOGIC_X1Y176_O = RIOB33_X105Y175_IOB_X1Y176_I;
  assign RIOI3_X105Y175_ILOGIC_X1Y175_O = RIOB33_X105Y175_IOB_X1Y175_I;
  assign RIOI3_X105Y177_ILOGIC_X1Y178_O = RIOB33_X105Y177_IOB_X1Y178_I;
  assign RIOI3_X105Y177_ILOGIC_X1Y177_O = RIOB33_X105Y177_IOB_X1Y177_I;
  assign RIOI3_X105Y179_ILOGIC_X1Y180_O = RIOB33_X105Y179_IOB_X1Y180_I;
  assign RIOI3_X105Y179_ILOGIC_X1Y179_O = RIOB33_X105Y179_IOB_X1Y179_I;
  assign RIOI3_X105Y183_ILOGIC_X1Y184_O = RIOB33_X105Y183_IOB_X1Y184_I;
  assign RIOI3_X105Y183_ILOGIC_X1Y183_O = RIOB33_X105Y183_IOB_X1Y183_I;
  assign RIOI3_X105Y185_ILOGIC_X1Y186_O = RIOB33_X105Y185_IOB_X1Y186_I;
  assign RIOI3_X105Y185_ILOGIC_X1Y185_O = RIOB33_X105Y185_IOB_X1Y185_I;
  assign RIOI3_X105Y189_ILOGIC_X1Y190_O = RIOB33_X105Y189_IOB_X1Y190_I;
  assign RIOI3_X105Y189_ILOGIC_X1Y189_O = RIOB33_X105Y189_IOB_X1Y189_I;
  assign RIOI3_X105Y191_ILOGIC_X1Y192_O = RIOB33_X105Y191_IOB_X1Y192_I;
  assign RIOI3_X105Y191_ILOGIC_X1Y191_O = RIOB33_X105Y191_IOB_X1Y191_I;
  assign RIOI3_X105Y195_ILOGIC_X1Y196_O = RIOB33_X105Y195_IOB_X1Y196_I;
  assign RIOI3_X105Y195_ILOGIC_X1Y195_O = RIOB33_X105Y195_IOB_X1Y195_I;
  assign RIOI3_X105Y197_ILOGIC_X1Y198_O = RIOB33_X105Y197_IOB_X1Y198_I;
  assign RIOI3_X105Y197_ILOGIC_X1Y197_O = RIOB33_X105Y197_IOB_X1Y197_I;
  assign RIOI3_SING_X105Y50_ILOGIC_X1Y50_O = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign RIOI3_SING_X105Y99_ILOGIC_X1Y99_O = RIOB33_SING_X105Y99_IOB_X1Y99_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_ILOGIC_X1Y150_O = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOI3_SING_X105Y199_ILOGIC_X1Y199_O = RIOB33_SING_X105Y199_IOB_X1Y199_I;
  assign RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y58_O = RIOB33_X105Y57_IOB_X1Y58_I;
  assign RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y57_O = RIOB33_X105Y57_IOB_X1Y57_I;
  assign RIOI3_TBYTESRC_X105Y69_ILOGIC_X1Y70_O = RIOB33_X105Y69_IOB_X1Y70_I;
  assign RIOI3_TBYTESRC_X105Y69_ILOGIC_X1Y69_O = RIOB33_X105Y69_IOB_X1Y69_I;
  assign RIOI3_TBYTESRC_X105Y81_ILOGIC_X1Y82_O = RIOB33_X105Y81_IOB_X1Y82_I;
  assign RIOI3_TBYTESRC_X105Y81_ILOGIC_X1Y81_O = RIOB33_X105Y81_IOB_X1Y81_I;
  assign RIOI3_TBYTESRC_X105Y93_ILOGIC_X1Y94_O = RIOB33_X105Y93_IOB_X1Y94_I;
  assign RIOI3_TBYTESRC_X105Y93_ILOGIC_X1Y93_O = RIOB33_X105Y93_IOB_X1Y93_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_O = RIOB33_X105Y157_IOB_X1Y158_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_O = RIOB33_X105Y157_IOB_X1Y157_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_O = RIOB33_X105Y169_IOB_X1Y170_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_O = RIOB33_X105Y169_IOB_X1Y169_I;
  assign RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y182_O = RIOB33_X105Y181_IOB_X1Y182_I;
  assign RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y181_O = RIOB33_X105Y181_IOB_X1Y181_I;
  assign RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y194_O = RIOB33_X105Y193_IOB_X1Y194_I;
  assign RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y193_O = RIOB33_X105Y193_IOB_X1Y193_I;
  assign RIOI3_TBYTETERM_X105Y63_ILOGIC_X1Y64_O = RIOB33_X105Y63_IOB_X1Y64_I;
  assign RIOI3_TBYTETERM_X105Y63_ILOGIC_X1Y63_O = RIOB33_X105Y63_IOB_X1Y63_I;
  assign RIOI3_TBYTETERM_X105Y87_ILOGIC_X1Y88_O = RIOB33_X105Y87_IOB_X1Y88_I;
  assign RIOI3_TBYTETERM_X105Y87_ILOGIC_X1Y87_O = RIOB33_X105Y87_IOB_X1Y87_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y164_O = RIOB33_X105Y163_IOB_X1Y164_I;
  assign RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_O = RIOB33_X105Y163_IOB_X1Y163_I;
  assign RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y188_O = RIOB33_X105Y187_IOB_X1Y188_I;
  assign RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y187_O = RIOB33_X105Y187_IOB_X1Y187_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D6 = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_A2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_A3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_A4 = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_A5 = RIOB33_X105Y53_IOB_X1Y53_I;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_A6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign LIOI3_SING_X0Y150_ILOGIC_X0Y150_D = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_B1 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_B2 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_B3 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_B4 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_B5 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_B6 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_C1 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_C2 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_C3 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_C4 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_C5 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_C6 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_D1 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_D2 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_D3 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_D4 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_D5 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X118Y115_D6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A4 = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A5 = CLBLL_L_X2Y123_SLICE_X0Y123_BQ;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_A1 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_A2 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_A3 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_A4 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_A5 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_A6 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_D1 = CLBLM_L_X70Y124_SLICE_X104Y124_AO6;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_B1 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_B2 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_B3 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_B4 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_B5 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_B6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B2 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y96_T1 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_C1 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_C2 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_C3 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_C4 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_C5 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_C6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B4 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_D1 = CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B5 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_D1 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_D2 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_D3 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_D4 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_D5 = 1'b1;
  assign CLBLL_R_X77Y115_SLICE_X119Y115_D6 = 1'b1;
  assign LIOI3_X0Y95_OLOGIC_X0Y95_T1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C2 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C6 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign LIOI3_X0Y155_ILOGIC_X0Y156_D = LIOB33_X0Y155_IOB_X0Y156_I;
  assign LIOI3_X0Y155_ILOGIC_X0Y155_D = LIOB33_X0Y155_IOB_X0Y155_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D6 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign RIOI3_X105Y77_ILOGIC_X1Y78_D = RIOB33_X105Y77_IOB_X1Y78_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_A1 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_A2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_A3 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_A6 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign RIOI3_X105Y77_ILOGIC_X1Y77_D = RIOB33_X105Y77_IOB_X1Y77_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_B1 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_B2 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_B3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_B4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_B6 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_C2 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_C3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_C4 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_C6 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y182_D = RIOB33_X105Y181_IOB_X1Y182_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign RIOI3_TBYTESRC_X105Y181_ILOGIC_X1Y181_D = RIOB33_X105Y181_IOB_X1Y181_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_D1 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_D2 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_D3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_D4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_D5 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X74Y115_SLICE_X113Y115_D6 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_A1 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_A2 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_A3 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_A4 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_A5 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_A6 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_B1 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_B2 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_B3 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_B4 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_B5 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_B6 = 1'b1;
  assign LIOI3_SING_X0Y199_ILOGIC_X0Y199_D = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_C1 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_C2 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_C3 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_C4 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_C5 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_C6 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_D1 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_D2 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_D3 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_D4 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_D5 = 1'b1;
  assign CLBLM_L_X74Y115_SLICE_X112Y115_D6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B4 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B5 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B6 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C4 = CLBLL_R_X73Y126_SLICE_X111Y126_F7AMUX_O;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C5 = CLBLM_R_X59Y117_SLICE_X88Y117_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_AX = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A1 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A2 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A3 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A4 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A5 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_A6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B1 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B2 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B3 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B4 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B5 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_B6 = 1'b1;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_A2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_A3 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_A4 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_A5 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_A6 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C1 = 1'b1;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C2 = 1'b1;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_B1 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_B2 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C4 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C5 = 1'b1;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_C1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_C2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_C3 = CLBLM_L_X70Y121_SLICE_X104Y121_DO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_C4 = CLBLM_L_X74Y116_SLICE_X113Y116_F7AMUX_O;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_C5 = CLBLM_L_X74Y115_SLICE_X113Y115_F8MUX_O;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_C6 = CLBLL_R_X75Y116_SLICE_X115Y116_F7AMUX_O;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D1 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D2 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D3 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D4 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D5 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_D6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A1 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A2 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_D1 = 1'b1;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_D2 = 1'b1;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_D3 = 1'b1;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_D4 = 1'b1;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_D5 = 1'b1;
  assign CLBLM_L_X74Y116_SLICE_X113Y116_D6 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A4 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_A6 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B1 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_A1 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_A2 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_A4 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_A6 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B4 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B5 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_B2 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_B3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_B4 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_B5 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C3 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C4 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C5 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_C1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_C2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_C4 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_C5 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_C6 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D2 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D3 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D4 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D5 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y61_ILOGIC_X1Y62_D = RIOB33_X105Y61_IOB_X1Y62_I;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_D1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_D2 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_D3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_D4 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_D5 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLM_L_X74Y116_SLICE_X112Y116_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_SING_X0Y200_ILOGIC_X0Y200_D = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLM_L_X56Y116_SLICE_X84Y116_AO6;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign RIOI3_X105Y61_ILOGIC_X1Y61_D = RIOB33_X105Y61_IOB_X1Y61_I;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_D1 = CLBLL_R_X71Y131_SLICE_X106Y131_AO6;
  assign LIOI3_X0Y97_OLOGIC_X0Y98_T1 = 1'b1;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_D1 = CLBLM_L_X70Y124_SLICE_X104Y124_CO6;
  assign LIOI3_X0Y97_OLOGIC_X0Y97_T1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B4 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A2 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A3 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A4 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A5 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B2 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B3 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B4 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_B6 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A3 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A5 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_A6 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C2 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B1 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B2 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B4 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_B6 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C5 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C2 = CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C3 = CLBLM_L_X74Y117_SLICE_X112Y117_F8MUX_O;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C4 = CLBLM_L_X74Y117_SLICE_X113Y117_F7AMUX_O;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_C6 = CLBLL_R_X75Y117_SLICE_X114Y117_F7AMUX_O;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D1 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D2 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D4 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_D6 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A2 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D2 = CLBLM_L_X74Y118_SLICE_X113Y118_F7AMUX_O;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D4 = CLBLL_R_X75Y117_SLICE_X115Y117_F8MUX_O;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D5 = CLBLM_L_X70Y121_SLICE_X104Y121_DO6;
  assign CLBLM_L_X74Y117_SLICE_X113Y117_D6 = CLBLL_R_X75Y117_SLICE_X114Y117_F7BMUX_O;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A5 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_A6 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A2 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A3 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A4 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_A6 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B4 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B5 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B3 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B4 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B5 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_B6 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C6 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C5 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C2 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C3 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C4 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_C6 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D2 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D4 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D5 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_D6 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D1 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D3 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D4 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y117_SLICE_X112Y117_D6 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y79_ILOGIC_X1Y80_D = RIOB33_X105Y79_IOB_X1Y80_I;
  assign RIOI3_X105Y79_ILOGIC_X1Y79_D = RIOB33_X105Y79_IOB_X1Y79_I;
  assign RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y194_D = RIOB33_X105Y193_IOB_X1Y194_I;
  assign RIOI3_TBYTESRC_X105Y193_ILOGIC_X1Y193_D = RIOB33_X105Y193_IOB_X1Y193_I;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C6 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A2 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A4 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A5 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_A6 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B2 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B4 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B5 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_B6 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C3 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_C6 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D3 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X113Y118_D6 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A3 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_A6 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B3 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_B6 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C3 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_C6 = 1'b1;
  assign LIOI3_X0Y159_ILOGIC_X0Y160_D = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D1 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D2 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D3 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D4 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D5 = 1'b1;
  assign CLBLM_L_X74Y118_SLICE_X112Y118_D6 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_A1 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_A2 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_A3 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_A4 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_A5 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_A6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A3 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_B1 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_B2 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_B3 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_B4 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_B5 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_B6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A6 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_C1 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_C2 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_C3 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_C4 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_C5 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_C6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C2 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_D1 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_D2 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_D3 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_D4 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_D5 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X71Y116_D6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D5 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_A1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_A2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_A4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_A5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_A6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_B1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_B2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_B3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_B6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A6 = CLBLL_R_X71Y125_SLICE_X106Y125_DO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B1 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_C1 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_C2 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_C3 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_C4 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_C5 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_C6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C5 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_D1 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_D2 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_D3 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_D4 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_D5 = 1'b1;
  assign CLBLM_L_X46Y116_SLICE_X70Y116_D6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D1 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D5 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_D6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A1 = CLBLM_L_X72Y131_SLICE_X108Y131_DO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A3 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A4 = CLBLM_L_X72Y131_SLICE_X108Y131_BO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_A6 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_AX = CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A4 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A5 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_A6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B2 = CLBLL_R_X71Y131_SLICE_X107Y131_CQ;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B4 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B5 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A1 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A2 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A5 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_A6 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B5 = RIOB33_X105Y169_IOB_X1Y170_I;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B1 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B2 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_B6 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B3 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_B6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C5 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C1 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C2 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C4 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_C6 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D3 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D4 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D5 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_D6 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D1 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D2 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D4 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y119_SLICE_X113Y119_D6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C1 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A4 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A6 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C2 = CLBLM_L_X72Y128_SLICE_X109Y128_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A1 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A2 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A4 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C3 = CLBLM_L_X74Y128_SLICE_X112Y128_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_A6 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B4 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B5 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C4 = CLBLL_R_X73Y129_SLICE_X110Y129_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B1 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C5 = CLBLM_L_X72Y128_SLICE_X109Y128_DO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_B6 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_C6 = CLBLL_R_X75Y127_SLICE_X114Y127_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C2 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C3 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C5 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_C6 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D2 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D3 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D4 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D5 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_D6 = 1'b1;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D2 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D3 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y119_SLICE_X112Y119_D6 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D4 = CLBLL_R_X73Y129_SLICE_X110Y129_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D1 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D5 = CLBLM_L_X72Y128_SLICE_X109Y128_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A2 = CLBLL_R_X71Y125_SLICE_X106Y125_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A4 = CLBLL_L_X2Y123_SLICE_X1Y123_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A6 = CLBLL_L_X2Y124_SLICE_X0Y124_AQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C6 = 1'b1;
  assign LIOI3_X0Y161_ILOGIC_X0Y162_D = LIOB33_X0Y161_IOB_X0Y162_I;
  assign LIOI3_X0Y161_ILOGIC_X0Y161_D = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D3 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D6 = 1'b1;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C2 = 1'b1;
  assign RIOI3_X105Y83_ILOGIC_X1Y84_D = RIOB33_X105Y83_IOB_X1Y84_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign RIOI3_X105Y83_ILOGIC_X1Y83_D = RIOB33_X105Y83_IOB_X1Y83_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C4 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C5 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C6 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B2 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A1 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A2 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A3 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A4 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A5 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_A6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B1 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B2 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B3 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B4 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B5 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_B6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A1 = CLBLM_L_X74Y121_SLICE_X113Y121_F8MUX_O;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A3 = CLBLM_L_X74Y119_SLICE_X113Y119_F7BMUX_O;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A4 = CLBLM_L_X74Y119_SLICE_X113Y119_F7AMUX_O;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_A6 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C1 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C2 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B1 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B2 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_A1 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_A2 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_A3 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_A4 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_A6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B3 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B4 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B5 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_B1 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_B2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_B4 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_B5 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_B6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C1 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C2 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C3 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_C2 = CLBLM_L_X72Y115_SLICE_X109Y115_F7BMUX_O;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_C3 = CLBLL_R_X71Y119_SLICE_X106Y119_AO6;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_C4 = CLBLM_L_X72Y114_SLICE_X109Y114_F7AMUX_O;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_C5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_C6 = CLBLL_R_X73Y114_SLICE_X110Y114_F8MUX_O;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D1 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D2 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D3 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D4 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D5 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_D6 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_D1 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_D2 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_D3 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_D4 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_D5 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X109Y114_D6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A2 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A3 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A4 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_A6 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_A1 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_A2 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_A3 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_A4 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_A5 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_A6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B2 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B3 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_B1 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_B2 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_B3 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_B4 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_B5 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_B6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C2 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C3 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_C1 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_C2 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_C3 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_C4 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_C5 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_C6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D1 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D2 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D3 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_D6 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_D1 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_D2 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_D3 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_D4 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_D5 = 1'b1;
  assign CLBLM_L_X72Y114_SLICE_X108Y114_D6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B2 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B5 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C4 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C5 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A2 = RIOB33_X105Y89_IOB_X1Y89_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A5 = LIOB33_X0Y195_IOB_X0Y195_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_A6 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C3 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B4 = LIOB33_X0Y177_IOB_X0Y178_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B5 = RIOB33_X105Y71_IOB_X1Y72_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C5 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C1 = RIOB33_X105Y195_IOB_X1Y196_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C4 = RIOB33_X105Y95_IOB_X1Y96_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_C6 = LIOB33_X0Y201_IOB_X0Y202_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A1 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A2 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A3 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A5 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_A6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D4 = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_A1 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_A2 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_A4 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_A6 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D5 = RIOB33_X105Y189_IOB_X1Y189_I;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X77Y122_SLICE_X118Y122_D6 = RIOB33_X105Y73_IOB_X1Y73_I;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_B1 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_B2 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_B5 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_B6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C1 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C2 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_C2 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_C3 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_C4 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_C5 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_C6 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D1 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D2 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A1 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A2 = 1'b1;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A3 = 1'b1;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_D1 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_D2 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_D4 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_D5 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X72Y115_SLICE_X109Y115_D6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A4 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A5 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B3 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B5 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B1 = 1'b1;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_A1 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_A2 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_A3 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_A4 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_A6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C2 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C3 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C4 = 1'b1;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C5 = 1'b1;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_B1 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_B2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_B3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_B6 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C6 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D2 = 1'b1;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D3 = 1'b1;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_C1 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_C2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D4 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D5 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D6 = 1'b1;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_C3 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_C4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_C6 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D2 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D3 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_D1 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_D2 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_D3 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_D4 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y115_SLICE_X108Y115_D6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A2 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A3 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A4 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A5 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_D1 = CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y88_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_D1 = CLBLL_R_X71Y119_SLICE_X106Y119_AO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B2 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y87_OLOGIC_X0Y87_T1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B3 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B5 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_B6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C2 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C3 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C5 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_C6 = 1'b1;
  assign LIOI3_X0Y165_ILOGIC_X0Y166_D = LIOB33_X0Y165_IOB_X0Y166_I;
  assign LIOI3_X0Y165_ILOGIC_X0Y165_D = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D2 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D3 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D5 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A1 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A2 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A4 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_A6 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X76Y133_SLICE_X116Y133_D6 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B2 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B5 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_B6 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign RIOI3_X105Y85_ILOGIC_X1Y86_D = RIOB33_X105Y85_IOB_X1Y86_I;
  assign RIOI3_X105Y85_ILOGIC_X1Y85_D = RIOB33_X105Y85_IOB_X1Y85_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C1 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C2 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_C6 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D1 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D3 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D5 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X72Y116_SLICE_X109Y116_D6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A1 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A4 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_A6 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B1 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B2 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_B6 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C1 = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C2 = CLBLM_L_X72Y116_SLICE_X109Y116_F7AMUX_O;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C4 = CLBLM_L_X72Y117_SLICE_X108Y117_F7AMUX_O;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C5 = CLBLM_L_X74Y116_SLICE_X112Y116_F8MUX_O;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_C6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D1 = CLBLM_L_X72Y117_SLICE_X108Y117_F7BMUX_O;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D2 = CLBLM_L_X70Y124_SLICE_X104Y124_CO6;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D3 = CLBLM_L_X72Y115_SLICE_X108Y115_F8MUX_O;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D4 = CLBLM_L_X72Y116_SLICE_X108Y116_F7AMUX_O;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y116_SLICE_X108Y116_D6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y58_D = RIOB33_X105Y57_IOB_X1Y58_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_L_X70Y123_SLICE_X105Y123_AO6;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_A1 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_A2 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_A3 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_A4 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_A5 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_A6 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_B1 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_B2 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_B3 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_B4 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_B5 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_B6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A4 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A5 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_A6 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_C1 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_C2 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B2 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A1 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A5 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_A6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B3 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B5 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B1 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B2 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B5 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_B6 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C1 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C2 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C2 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C3 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C4 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C5 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_C6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D1 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D2 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D3 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D5 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_D6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D1 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D2 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D3 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D4 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D5 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X109Y117_D6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_A6 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A1 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A4 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A5 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_A6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B2 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B3 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B1 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B2 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B4 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_B6 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C1 = CLBLM_L_X74Y124_SLICE_X113Y124_F7BMUX_O;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C2 = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C3 = CLBLM_L_X74Y123_SLICE_X113Y123_F8MUX_O;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C1 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C4 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C5 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_C6 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D4 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D5 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D1 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D2 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_D3 = 1'b1;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLM_L_X70Y123_SLICE_X104Y123_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D1 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D2 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X72Y117_SLICE_X108Y117_D6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A5 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A6 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_A1 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_A2 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_A3 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_A4 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_A5 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_A6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_B1 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_B2 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_B3 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_B4 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_B5 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_B6 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_C1 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_C2 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_C3 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_C4 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_C5 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_C6 = 1'b1;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_D3 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_D1 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_D2 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_D3 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_D4 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_D5 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X89Y117_D6 = 1'b1;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_D5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_A1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_A2 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_A3 = CLBLM_R_X59Y117_SLICE_X88Y117_AQ;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_A4 = CLBLM_R_X59Y118_SLICE_X88Y118_AQ;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_A5 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_A6 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_AX = CLBLM_R_X59Y118_SLICE_X88Y118_AO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_B1 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_B2 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_B3 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_B4 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_B5 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_B6 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_C1 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_C2 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_C3 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_C4 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_C5 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_C6 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLM_L_X56Y116_SLICE_X84Y116_AO6;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign RIOI3_SING_X105Y50_ILOGIC_X1Y50_D = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_D1 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_D2 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_D3 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_D4 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_D5 = 1'b1;
  assign CLBLM_R_X59Y117_SLICE_X88Y117_D6 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_L_X70Y122_SLICE_X104Y122_AO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y183_ILOGIC_X1Y184_D = RIOB33_X105Y183_IOB_X1Y184_I;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A3 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_A6 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B2 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B3 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B4 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B5 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign RIOI3_X105Y183_ILOGIC_X1Y183_D = RIOB33_X105Y183_IOB_X1Y183_I;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C1 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C2 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C3 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C4 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_C6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D5 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_D2 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D1 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D2 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D4 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D5 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X77Y125_SLICE_X118Y125_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_A2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_A3 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_A4 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_A6 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_B1 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_B2 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A1 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A2 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A4 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_A6 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_B3 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_B5 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B2 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B3 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_B6 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A2 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A4 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A5 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_A6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C2 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B2 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B4 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B5 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_B6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C2 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D4 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D5 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D6 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C4 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C5 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_C6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A1 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A2 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D1 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D2 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D3 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D4 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D5 = 1'b1;
  assign CLBLL_R_X77Y125_SLICE_X119Y125_D6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A4 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B1 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B2 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B3 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B5 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_B6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_C1 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_C3 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C2 = CLBLM_L_X72Y118_SLICE_X109Y118_F7AMUX_O;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C4 = CLBLM_L_X72Y117_SLICE_X109Y117_F7AMUX_O;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C5 = CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_C6 = CLBLL_R_X71Y118_SLICE_X107Y118_F8MUX_O;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_D1 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_D2 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_D3 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_D4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_D6 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign LIOI3_X0Y167_ILOGIC_X0Y168_D = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D2 = CLBLL_R_X73Y118_SLICE_X110Y118_F8MUX_O;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D3 = CLBLM_L_X72Y118_SLICE_X109Y118_F7BMUX_O;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D4 = CLBLM_L_X72Y118_SLICE_X108Y118_F7AMUX_O;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D5 = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_D6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign LIOI3_X0Y167_ILOGIC_X0Y167_D = LIOB33_X0Y167_IOB_X0Y167_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y152_D = RIOB33_X105Y151_IOB_X1Y152_I;
  assign RIOI3_X105Y151_ILOGIC_X1Y151_D = RIOB33_X105Y151_IOB_X1Y151_I;
  assign RIOI3_X105Y89_ILOGIC_X1Y90_D = RIOB33_X105Y89_IOB_X1Y90_I;
  assign RIOI3_X105Y89_ILOGIC_X1Y89_D = RIOB33_X105Y89_IOB_X1Y89_I;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_A1 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_A2 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_A3 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_A4 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_A5 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_A6 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_B1 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_B2 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_B3 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_B4 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_B5 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_B6 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_C1 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_C2 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_C3 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_C4 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_C5 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_C6 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_D1 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_D2 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_D3 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_D4 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_D5 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X89Y118_D6 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_A1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_A2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_A3 = CLBLM_R_X59Y118_SLICE_X88Y118_AQ;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_A4 = CLBLM_R_X59Y118_SLICE_X88Y118_BO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_A5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_A6 = CLBLL_R_X73Y122_SLICE_X110Y122_BO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B6 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_AX = CLBLM_R_X59Y117_SLICE_X88Y117_AO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_B2 = RIOB33_X105Y163_IOB_X1Y164_I;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_B3 = CLBLM_R_X59Y118_SLICE_X88Y118_AQ;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_B4 = CLBLM_R_X59Y117_SLICE_X88Y117_AQ;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_B6 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_C1 = 1'b1;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_D3 = CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_C2 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_C3 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_C4 = 1'b1;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_D4 = CLBLM_L_X72Y119_SLICE_X108Y119_CO6;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_C5 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_C6 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_D1 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_D2 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_D3 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_D4 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_D5 = 1'b1;
  assign CLBLM_R_X59Y118_SLICE_X88Y118_D6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C4 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A3 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C5 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C6 = 1'b1;
  assign RIOI3_SING_X105Y99_ILOGIC_X1Y99_D = RIOB33_SING_X105Y99_IOB_X1Y99_I;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B2 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A2 = LIOB33_X0Y189_IOB_X0Y190_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A3 = RIOB33_X105Y83_IOB_X1Y84_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A4 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_A6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B1 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B2 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B3 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B4 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B5 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_B6 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A1 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A2 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A5 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C1 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_C2 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B2 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A1 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A2 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A5 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_A6 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B3 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B4 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_B5 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B1 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B3 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B4 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C2 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_B6 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_C1 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C3 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C1 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C2 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C3 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C4 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D1 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C5 = 1'b1;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D2 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y125_SLICE_X113Y125_D4 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C6 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D1 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D2 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D3 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D4 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y119_SLICE_X109Y119_D6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A1 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A2 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_A6 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A1 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A2 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A5 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_A6 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B1 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B1 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B5 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_B6 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C1 = CLBLM_L_X74Y126_SLICE_X112Y126_F8MUX_O;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C2 = CLBLM_L_X74Y125_SLICE_X113Y125_F7AMUX_O;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_C3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C2 = CLBLM_L_X72Y119_SLICE_X109Y119_F7AMUX_O;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C3 = CLBLL_R_X73Y119_SLICE_X110Y119_F8MUX_O;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C4 = CLBLM_L_X72Y119_SLICE_X108Y119_F7AMUX_O;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C5 = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D2 = CLBLM_L_X74Y125_SLICE_X113Y125_F7BMUX_O;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D4 = CLBLM_L_X74Y124_SLICE_X113Y124_F7AMUX_O;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D5 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLM_L_X74Y125_SLICE_X112Y125_D6 = CLBLL_R_X73Y125_SLICE_X111Y125_F8MUX_O;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D1 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D2 = CLBLM_L_X72Y119_SLICE_X109Y119_F7BMUX_O;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D3 = CLBLL_R_X71Y119_SLICE_X107Y119_F7AMUX_O;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D2 = 1'b1;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D5 = CLBLM_L_X72Y121_SLICE_X108Y121_F8MUX_O;
  assign CLBLM_L_X72Y119_SLICE_X108Y119_D6 = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D4 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B4 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B6 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_C2 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_C3 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_C5 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_C6 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C4 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A1 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A2 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A3 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A4 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A5 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_A6 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B1 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B2 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A2 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A3 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_A6 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B3 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B4 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_B5 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B1 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B2 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B4 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B5 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_B4 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C1 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_C3 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C1 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C2 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C3 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_C6 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D1 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D2 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D3 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D4 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y126_SLICE_X113Y126_D5 = 1'b1;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D2 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D5 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X72Y120_SLICE_X109Y120_D6 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D4 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A1 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A2 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D5 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A3 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A1 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A2 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A3 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A4 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D6 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_C1 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B1 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_B3 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B1 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B2 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B3 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B4 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_C2 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C1 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_C3 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C1 = CLBLL_R_X71Y122_SLICE_X106Y122_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C2 = CLBLM_L_X74Y120_SLICE_X113Y120_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C3 = CLBLL_R_X71Y120_SLICE_X107Y120_AO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C4 = CLBLL_R_X73Y120_SLICE_X111Y120_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C5 = CLBLM_L_X72Y120_SLICE_X108Y120_DO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_C6 = CLBLL_R_X73Y120_SLICE_X111Y120_CO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D1 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D2 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D3 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D5 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_D6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D2 = CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D4 = CLBLM_L_X72Y120_SLICE_X108Y120_F7AMUX_O;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D5 = CLBLM_L_X72Y121_SLICE_X109Y121_F8MUX_O;
  assign CLBLM_L_X72Y120_SLICE_X108Y120_D6 = CLBLL_R_X71Y120_SLICE_X106Y120_F7BMUX_O;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_A1 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_A2 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_A3 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_A4 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_A5 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_A6 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_B1 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_B2 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_B3 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_B4 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_B5 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_B6 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_C1 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_C2 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_C3 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_C4 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_C5 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_C6 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_D1 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_D2 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_D3 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_D4 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_D5 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X67Y118_D6 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_A1 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_A2 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_A4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_A5 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_A6 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_B1 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_B2 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_B3 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_B4 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_B5 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_B6 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_C1 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_C2 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_C3 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_C4 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_C5 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_C6 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_D1 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_D2 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_D3 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_D4 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_D5 = 1'b1;
  assign CLBLM_L_X44Y118_SLICE_X66Y118_D6 = 1'b1;
  assign LIOI3_X0Y171_ILOGIC_X0Y172_D = LIOB33_X0Y171_IOB_X0Y172_I;
  assign LIOI3_X0Y171_ILOGIC_X0Y171_D = LIOB33_X0Y171_IOB_X0Y171_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y154_D = RIOB33_X105Y153_IOB_X1Y154_I;
  assign RIOI3_X105Y153_ILOGIC_X1Y153_D = RIOB33_X105Y153_IOB_X1Y153_I;
  assign RIOI3_X105Y91_ILOGIC_X1Y92_D = RIOB33_X105Y91_IOB_X1Y92_I;
  assign RIOI3_X105Y91_ILOGIC_X1Y91_D = RIOB33_X105Y91_IOB_X1Y91_I;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A2 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A3 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A4 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_A6 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B1 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A2 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A3 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A4 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_A6 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B2 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B3 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B4 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B5 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C1 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C2 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_C3 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C1 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C3 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C4 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_C6 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D1 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D2 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D3 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D4 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D5 = 1'b1;
  assign CLBLM_L_X74Y127_SLICE_X113Y127_D6 = 1'b1;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D1 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D4 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D5 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X72Y121_SLICE_X109Y121_D6 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A1 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A4 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_A6 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A1 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A3 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A4 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A5 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B1 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B2 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_B3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B1 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B3 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B4 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_B6 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C2 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_C3 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C2 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C3 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_C6 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D2 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D3 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D4 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D5 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X74Y127_SLICE_X112Y127_D6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D2 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D3 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D5 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X72Y121_SLICE_X108Y121_D6 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C3 = 1'b1;
  assign CLBLM_L_X76Y124_SLICE_X117Y124_C6 = 1'b1;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A3 = RIOB33_X105Y69_IOB_X1Y69_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A5 = LIOB33_X0Y175_IOB_X0Y175_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_A6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B2 = LIOB33_X0Y201_IOB_X0Y201_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B3 = RIOB33_X105Y195_IOB_X1Y195_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B5 = RIOB33_X105Y95_IOB_X1Y95_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_B6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C2 = LIOB33_X0Y193_IOB_X0Y194_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C5 = RIOB33_X105Y87_IOB_X1Y88_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_C6 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D1 = LIOB33_SING_X0Y200_IOB_X0Y200_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D3 = RIOB33_X105Y193_IOB_X1Y194_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D5 = RIOB33_X105Y93_IOB_X1Y94_I;
  assign CLBLL_R_X77Y129_SLICE_X118Y129_D6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A1 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A5 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A1 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A2 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A3 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A4 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A5 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_A6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A1 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A4 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A5 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_A2 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B4 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B5 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B1 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B3 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B4 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B5 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_B6 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_A3 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C3 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C4 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C5 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_C1 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_B2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_B3 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_B4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_B6 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_C1 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_C2 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_C3 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_C4 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_C5 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D3 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_C6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D5 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X109Y122_D6 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D2 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D3 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D5 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D6 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_D1 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_D2 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_D3 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_D4 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_D5 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_D6 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A1 = CLBLM_L_X72Y123_SLICE_X109Y123_F8MUX_O;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A2 = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A4 = CLBLM_L_X72Y123_SLICE_X108Y123_F7BMUX_O;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_A6 = CLBLM_L_X72Y123_SLICE_X108Y123_F7AMUX_O;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B1 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B2 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B3 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B4 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B5 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_B6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C3 = CLBLL_R_X75Y128_SLICE_X114Y128_F8MUX_O;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C1 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C2 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C3 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C4 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C5 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_C6 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_A1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_A3 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_A4 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_A5 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_A6 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D1 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D2 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_B1 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_B3 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_B4 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_B5 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_B6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D1 = 1'b1;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D2 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y122_SLICE_X108Y122_D3 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_C1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_C2 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_C3 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_C4 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_C6 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D2 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_D1 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_D2 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_D3 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_D4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y115_SLICE_X115Y115_D6 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D3 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_L_X72Y131_SLICE_X108Y131_AO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D4 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_C6 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D5 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B4 = RIOB33_X105Y151_IOB_X1Y152_I;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B6 = CLBLM_L_X70Y128_SLICE_X105Y128_AQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_BX = CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C1 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C2 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C3 = CLBLM_L_X70Y128_SLICE_X105Y128_BQ;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A1 = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A4 = RIOB33_X105Y193_IOB_X1Y193_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A5 = RIOB33_X105Y77_IOB_X1Y77_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_A6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C5 = CLBLM_L_X70Y128_SLICE_X105Y128_AQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B3 = RIOB33_X105Y187_IOB_X1Y188_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B5 = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_B6 = RIOB33_X105Y63_IOB_X1Y63_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C1 = LIOB33_X0Y203_IOB_X0Y203_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C3 = RIOB33_X105Y97_IOB_X1Y97_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C5 = RIOB33_X105Y197_IOB_X1Y197_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_C6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D3 = LIOB33_X0Y177_IOB_X0Y177_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D5 = RIOB33_X105Y71_IOB_X1Y71_I;
  assign CLBLL_R_X77Y130_SLICE_X118Y130_D6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A2 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A3 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A1 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A2 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A3 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A4 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A5 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_A6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A4 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A5 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_A1 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_A3 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B4 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B5 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B6 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_A5 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_A6 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B1 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B2 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_A1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C3 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C4 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C5 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C6 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_A2 = CLBLL_R_X71Y117_SLICE_X106Y117_F7AMUX_O;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_A3 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_A4 = CLBLL_R_X71Y117_SLICE_X106Y117_F7BMUX_O;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_A5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_A6 = CLBLL_R_X71Y116_SLICE_X106Y116_F8MUX_O;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_B1 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_B2 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_B3 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_B4 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_B5 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_B6 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_C2 = CLBLL_R_X75Y115_SLICE_X114Y115_F7AMUX_O;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_C1 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_C4 = CLBLL_R_X75Y116_SLICE_X114Y116_F7AMUX_O;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_C5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_C4 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D2 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D3 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D4 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D5 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D6 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_D1 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_D2 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_D3 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_D4 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_D5 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_D6 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_D1 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_D2 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_D3 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_D4 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_D5 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X105Y117_D6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A1 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A3 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A4 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A5 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_A1 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_A2 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_A3 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_A4 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_A5 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_A6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B2 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_A1 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_A2 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_A3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_B5 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_B6 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_A5 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_A6 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_B1 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_B2 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_B3 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_B1 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_C3 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_C4 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_C5 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_C6 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_B2 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_B3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_B5 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_C1 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_C2 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_C3 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_C4 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_C5 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_C6 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_D1 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_D2 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_D3 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_D4 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_D5 = 1'b1;
  assign CLBLM_L_X70Y117_SLICE_X104Y117_D6 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_D1 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_D2 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_D3 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_D4 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_D5 = 1'b1;
  assign CLBLL_R_X75Y116_SLICE_X115Y116_D6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B5 = CLBLM_L_X70Y127_SLICE_X104Y127_BQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A3 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign RIOI3_SING_X105Y199_ILOGIC_X1Y199_D = RIOB33_SING_X105Y199_IOB_X1Y199_I;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A4 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C3 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C4 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C5 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B2 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A5 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B4 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B5 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_B6 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C2 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A2 = LIOB33_X0Y197_IOB_X0Y197_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A3 = RIOB33_X105Y91_IOB_X1Y91_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A5 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_A6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C3 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C4 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B2 = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B3 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B4 = RIOB33_X105Y83_IOB_X1Y83_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B5 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_B6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A4 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C5 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C2 = LIOB33_X0Y195_IOB_X0Y196_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C5 = RIOB33_X105Y89_IOB_X1Y90_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_C6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A5 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_C6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D1 = RIOB33_X105Y69_IOB_X1Y70_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D2 = LIOB33_X0Y175_IOB_X0Y176_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D5 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y131_SLICE_X118Y131_D6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B2 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B3 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B4 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D1 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A1 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A2 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A3 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A4 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A5 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_A6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D2 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_A1 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_A2 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_A3 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B4 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B5 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A6 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C3 = 1'b1;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C5 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B3 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_B1 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_B2 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_B3 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_B4 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C1 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C1 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C2 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_C1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_C2 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_C3 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_C4 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_C6 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D2 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D3 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D4 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D5 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D6 = 1'b1;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_D1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_D2 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_D3 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_D4 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_D6 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C5 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C6 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D4 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D5 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A2 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A4 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A5 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_A6 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A1 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B1 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B4 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B5 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_B6 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A3 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_A1 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_A2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_A4 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_A5 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_A6 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C1 = CLBLM_L_X70Y123_SLICE_X104Y123_BO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C2 = CLBLM_L_X72Y124_SLICE_X109Y124_F7AMUX_O;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_B1 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_B2 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_B4 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_B6 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C4 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C5 = CLBLL_R_X73Y124_SLICE_X110Y124_F8MUX_O;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_C1 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_C2 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_C4 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_C6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D1 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D1 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D2 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D3 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D4 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D5 = 1'b1;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_D1 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_D2 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_D3 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_D4 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X115Y117_D6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B1 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D4 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D5 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B3 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_D6 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B4 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_B6 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C2 = CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C4 = CLBLM_L_X74Y128_SLICE_X112Y128_F7AMUX_O;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C5 = CLBLM_L_X74Y127_SLICE_X112Y127_F7BMUX_O;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_C6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B3 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X70Y121_SLICE_X105Y121_AO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D3 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D4 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_L_X70Y122_SLICE_X104Y122_CO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D5 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_D6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C1 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C2 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C5 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_C6 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_A2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_A3 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_A4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_A5 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_A6 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_B2 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_B3 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_B4 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_B6 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B2 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B4 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B5 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_B6 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_C2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C1 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C2 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_C4 = CLBLL_R_X75Y118_SLICE_X114Y118_F7AMUX_O;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C6 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A6 = CLBLL_R_X71Y116_SLICE_X107Y116_CO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_AX = CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_D1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_D2 = 1'b1;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_D3 = 1'b1;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_D4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_D5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D1 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D2 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D3 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D4 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C2 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C4 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C5 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C6 = RIOB33_X105Y177_IOB_X1Y177_I;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A2 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A4 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A5 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A6 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D2 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D3 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D4 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B1 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B2 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B3 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B5 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D5 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A1 = CLBLM_L_X70Y119_SLICE_X104Y119_BO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_A2 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C2 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C4 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C5 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_C6 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_B2 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_B3 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_B4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_B6 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_C1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_C2 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D4 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D6 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_C4 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_C5 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_C6 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C6 = CLBLM_L_X72Y118_SLICE_X108Y118_CO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_D1 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_D2 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_D3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_D4 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_D6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D2 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D5 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_D6 = 1'b1;
  assign LIOI3_X0Y175_ILOGIC_X0Y176_D = LIOB33_X0Y175_IOB_X0Y176_I;
  assign LIOI3_X0Y175_ILOGIC_X0Y175_D = LIOB33_X0Y175_IOB_X0Y175_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y160_D = RIOB33_X105Y159_IOB_X1Y160_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign RIOI3_X105Y159_ILOGIC_X1Y159_D = RIOB33_X105Y159_IOB_X1Y159_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign RIOI3_X105Y97_ILOGIC_X1Y98_D = RIOB33_X105Y97_IOB_X1Y98_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y188_D = LIOB33_X0Y187_IOB_X0Y188_I;
  assign RIOI3_X105Y97_ILOGIC_X1Y97_D = RIOB33_X105Y97_IOB_X1Y97_I;
  assign LIOI3_TBYTETERM_X0Y187_ILOGIC_X0Y187_D = LIOB33_X0Y187_IOB_X0Y187_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_A2 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_A3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_A4 = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_A5 = RIOB33_X105Y85_IOB_X1Y85_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_A6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_B1 = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_B2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_B3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_B4 = RIOB33_X105Y191_IOB_X1Y192_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_B5 = RIOB33_X105Y75_IOB_X1Y76_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_B6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_C1 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_C2 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_C3 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_C4 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_C5 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_C6 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_D1 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_D2 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_D3 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_D4 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_D5 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X118Y133_D6 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_A1 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_A2 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_A3 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_A4 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_A5 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_A6 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_A1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_A4 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_A5 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_A6 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_B1 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_B2 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_B3 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_B2 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_B3 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_B4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A1 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_B5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_B6 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B1 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B5 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_C2 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_C3 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_C4 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_C5 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_C6 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_D2 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_D3 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_D4 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_D5 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C6 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_D1 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_D2 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_D3 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_D4 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_D5 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_D6 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D1 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D4 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D5 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_D6 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A1 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A2 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A3 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A4 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_A2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_A3 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_A4 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_A5 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B4 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B5 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_A6 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B1 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C1 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C2 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C3 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_B1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C6 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_B2 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_B4 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_B5 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_B6 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_C1 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_C2 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_C3 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_C4 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_C5 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_C6 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D5 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D6 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_D1 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_D2 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_D3 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_D4 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_D5 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X115Y119_D6 = 1'b1;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C3 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X76Y125_SLICE_X117Y125_C6 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_B5 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_B6 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_A2 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_A3 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_A4 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_A5 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_A6 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_B2 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_B3 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_B4 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_B5 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A1 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_C1 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_C2 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_C4 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A6 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_C5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_C6 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A2 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B2 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B4 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B5 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_B6 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_A1 = CLBLM_L_X70Y121_SLICE_X105Y121_BO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_A3 = CLBLM_L_X70Y121_SLICE_X105Y121_AQ;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C2 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_D1 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C4 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C5 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_D2 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_D4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_D5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X75Y120_SLICE_X114Y120_D6 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_B2 = CLBLM_L_X70Y121_SLICE_X105Y121_BQ;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_B3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_B5 = RIOB33_X105Y173_IOB_X1Y174_I;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_B6 = CLBLM_L_X70Y121_SLICE_X105Y121_AQ;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_BX = CLBLM_L_X70Y121_SLICE_X105Y121_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D4 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D5 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_C1 = CLBLM_L_X70Y121_SLICE_X105Y121_BQ;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_C2 = RIOB33_X105Y175_IOB_X1Y175_I;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_C5 = CLBLM_L_X70Y121_SLICE_X105Y121_AQ;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_C6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A1 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A2 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A4 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_A6 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_D1 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_D3 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B1 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B2 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B3 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B4 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_A6 = CLBLL_R_X71Y119_SLICE_X106Y119_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_A1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C2 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C4 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C5 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_C6 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_C1 = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_C2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_C3 = CLBLM_L_X76Y120_SLICE_X116Y120_F8MUX_O;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_C4 = CLBLL_R_X75Y120_SLICE_X115Y120_F7AMUX_O;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_C5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_C1 = CLBLM_L_X70Y121_SLICE_X104Y121_BQ;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_C6 = CLBLL_R_X75Y119_SLICE_X115Y119_F7AMUX_O;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_C4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D2 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D4 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D5 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X72Y127_SLICE_X108Y127_D6 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_D1 = 1'b1;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_D2 = 1'b1;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_D3 = 1'b1;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_D4 = 1'b1;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_D5 = 1'b1;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_D6 = 1'b1;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_CX = CLBLM_L_X70Y121_SLICE_X104Y121_BO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_D1 = CLBLM_L_X70Y121_SLICE_X104Y121_BQ;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_D2 = CLBLM_L_X70Y121_SLICE_X104Y121_CQ;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_D3 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_D4 = RIOB33_X105Y179_IOB_X1Y179_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_D5 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_D6 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_DX = CLBLM_L_X70Y121_SLICE_X104Y121_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_B6 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C2 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X76Y125_SLICE_X116Y125_C3 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A4 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A5 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B2 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B3 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B4 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B5 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B6 = 1'b1;
  assign LIOI3_X0Y177_ILOGIC_X0Y178_D = LIOB33_X0Y177_IOB_X0Y178_I;
  assign LIOI3_X0Y177_ILOGIC_X0Y177_D = LIOB33_X0Y177_IOB_X0Y177_I;
  assign RIOI3_X105Y161_ILOGIC_X1Y162_D = RIOB33_X105Y161_IOB_X1Y162_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign RIOI3_X105Y161_ILOGIC_X1Y161_D = RIOB33_X105Y161_IOB_X1Y161_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y82_D = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_TBYTESRC_X0Y81_ILOGIC_X0Y81_D = LIOB33_X0Y81_IOB_X0Y81_I;
  assign RIOI3_TBYTETERM_X105Y63_ILOGIC_X1Y64_D = RIOB33_X105Y63_IOB_X1Y64_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_TBYTETERM_X105Y63_ILOGIC_X1Y63_D = RIOB33_X105Y63_IOB_X1Y63_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A1 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A4 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A5 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A6 = CLBLL_R_X71Y120_SLICE_X107Y120_CO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A1 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_AX = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B1 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B2 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B4 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A5 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_BX = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_A2 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_A3 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_A4 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_A5 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_A6 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_A1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C2 = CLBLL_R_X71Y116_SLICE_X107Y116_AO6;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_B1 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_B2 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_B3 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_B4 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_B5 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_B6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C6 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_CX = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_C1 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_C2 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_C3 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_C4 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_C5 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_C6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D3 = CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D5 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D6 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D3 = CLBLM_L_X74Y128_SLICE_X113Y128_F8MUX_O;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_D1 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_D2 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_D3 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_D4 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_D5 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X105Y122_D6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_A6 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_A1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_A3 = CLBLM_L_X70Y122_SLICE_X104Y122_AQ;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_A4 = CLBLM_L_X70Y122_SLICE_X104Y122_BO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_A6 = CLBLM_L_X70Y119_SLICE_X104Y119_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A6 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_AX = CLBLM_L_X70Y122_SLICE_X104Y122_CO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_B1 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_B2 = CLBLM_L_X70Y122_SLICE_X104Y122_BQ;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_B6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B3 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_BX = CLBLM_L_X70Y122_SLICE_X104Y122_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C6 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_C1 = CLBLM_L_X70Y122_SLICE_X104Y122_BQ;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_C2 = CLBLM_L_X70Y122_SLICE_X104Y122_AQ;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_C3 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_C5 = RIOB33_X105Y173_IOB_X1Y173_I;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_C6 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D6 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_D1 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_D2 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_D3 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_D4 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_D5 = 1'b1;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_D6 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_A1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_A6 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_A2 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_A3 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_A4 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_A5 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y164_D = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_B1 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_B2 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_B3 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_B4 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_B5 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_B6 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_A1 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_C1 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_C2 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_C3 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_A2 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_C4 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_C5 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B1 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_C6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B2 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_A4 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_D1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B3 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_D2 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_D4 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_D5 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B4 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_D6 = 1'b1;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X49Y116_SLICE_X75Y116_D3 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B5 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_A3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_B6 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_A4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_A5 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_A6 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y115_SLICE_X114Y115_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_B1 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_B2 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_B3 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_B4 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_B5 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_B6 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_C1 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_C2 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_C3 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_C4 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_C5 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_C6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C2 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_A1 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C3 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_D1 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_D2 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_D3 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_D4 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_D5 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C4 = 1'b1;
  assign CLBLM_R_X49Y116_SLICE_X74Y116_D6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C5 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_ILOGIC_X0Y163_D = LIOB33_X0Y163_IOB_X0Y163_I;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B2 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B4 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X74Y129_SLICE_X113Y129_D1 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_B6 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A1 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A1 = CLBLM_L_X70Y123_SLICE_X105Y123_AQ;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A4 = CLBLM_L_X70Y123_SLICE_X105Y123_BO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A5 = CLBLL_R_X73Y122_SLICE_X110Y122_CO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_A6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_AX = CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B1 = CLBLM_L_X70Y123_SLICE_X105Y123_AQ;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B2 = CLBLM_L_X70Y123_SLICE_X105Y123_BQ;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B5 = RIOB33_X105Y167_IOB_X1Y168_I;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_B6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_BX = CLBLM_L_X70Y123_SLICE_X105Y123_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C1 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C2 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C3 = CLBLM_L_X70Y123_SLICE_X105Y123_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C6 = RIOB33_X105Y169_IOB_X1Y169_I;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A1 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_C5 = CLBLM_L_X70Y123_SLICE_X105Y123_AQ;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C3 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_CX = CLBLM_L_X70Y123_SLICE_X105Y123_DO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C4 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A3 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D1 = CLBLM_L_X70Y124_SLICE_X105Y124_AO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D2 = CLBLM_L_X70Y124_SLICE_X105Y124_AQ;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D4 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D6 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A4 = CLBLM_L_X70Y119_SLICE_X105Y119_BO6;
  assign CLBLM_L_X70Y123_SLICE_X105Y123_D3 = CLBLL_R_X71Y120_SLICE_X107Y120_DO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_C6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A5 = CLBLM_L_X70Y121_SLICE_X104Y121_AQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A1 = CLBLM_L_X70Y121_SLICE_X104Y121_DQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A2 = RIOB33_X105Y165_IOB_X1Y166_I;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B2 = RIOB33_X105Y167_IOB_X1Y167_I;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B3 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B5 = CLBLM_L_X70Y121_SLICE_X104Y121_AQ;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C1 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C2 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B2 = CLBLM_L_X70Y119_SLICE_X105Y119_BQ;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = 1'b1;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B5 = RIOB33_X105Y175_IOB_X1Y176_I;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D2 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D4 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D5 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_B6 = CLBLM_L_X70Y119_SLICE_X105Y119_AQ;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D3 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B1 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B2 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B3 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_BX = CLBLM_L_X70Y119_SLICE_X105Y119_AO6;
  assign CLBLM_L_X72Y124_SLICE_X109Y124_D6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B4 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C1 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_L_X70Y127_SLICE_X104Y127_AO6;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_C3 = CLBLM_L_X70Y119_SLICE_X105Y119_BQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X70Y121_SLICE_X104Y121_DO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C2 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C3 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C4 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_D1 = CLBLM_L_X70Y129_SLICE_X104Y129_AO6;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y94_T1 = 1'b1;
  assign RIOI3_X105Y185_ILOGIC_X1Y186_D = RIOB33_X105Y185_IOB_X1Y186_I;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_D1 = CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  assign LIOI3_TBYTESRC_X0Y93_OLOGIC_X0Y93_T1 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D5 = 1'b1;
  assign RIOI3_X105Y185_ILOGIC_X1Y185_D = RIOB33_X105Y185_IOB_X1Y185_I;
  assign CLBLM_L_X70Y119_SLICE_X105Y119_D6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D1 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D2 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D3 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D4 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D5 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_D6 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A1 = CLBLL_R_X75Y124_SLICE_X114Y124_F8MUX_O;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A2 = CLBLM_L_X70Y121_SLICE_X105Y121_CO6;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A5 = CLBLL_R_X75Y124_SLICE_X115Y124_F7BMUX_O;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_A6 = CLBLL_R_X75Y124_SLICE_X115Y124_F7AMUX_O;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C3 = CLBLM_L_X72Y124_SLICE_X109Y124_F7BMUX_O;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B1 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B2 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A4 = CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B4 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B5 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_B6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C1 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C2 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C4 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C5 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_C6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_A6 = CLBLL_R_X71Y119_SLICE_X106Y119_CO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D1 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D2 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D4 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D5 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X114Y123_D6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A1 = RIOB33_X105Y181_IOB_X1Y182_I;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A2 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A3 = CLBLM_L_X70Y124_SLICE_X105Y124_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_A6 = CLBLM_L_X70Y123_SLICE_X105Y123_CQ;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_AX = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign LIOI3_X0Y179_ILOGIC_X0Y180_D = LIOB33_X0Y179_IOB_X0Y180_I;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B1 = RIOB33_X105Y183_IOB_X1Y183_I;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B2 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B2 = CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B3 = CLBLM_L_X70Y124_SLICE_X105Y124_AQ;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B5 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_B6 = CLBLM_L_X70Y123_SLICE_X105Y123_CQ;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B3 = CLBLM_L_X70Y119_SLICE_X104Y119_AQ;
  assign LIOI3_X0Y179_ILOGIC_X0Y179_D = LIOB33_X0Y179_IOB_X0Y179_I;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C1 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C2 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C3 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C4 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C5 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_C6 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A1 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A2 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A3 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_B6 = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_A4 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D1 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D2 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D3 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D4 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D5 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X105Y124_D6 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B1 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B2 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B4 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B5 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_B6 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C1 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C2 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C4 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C5 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_C6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A3 = CLBLM_L_X70Y124_SLICE_X104Y124_AQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A4 = CLBLM_L_X70Y124_SLICE_X104Y124_BO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A5 = CLBLL_R_X73Y122_SLICE_X110Y122_AO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C1 = CLBLM_L_X70Y117_SLICE_X105Y117_AO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B6 = CLBLM_L_X70Y124_SLICE_X104Y124_AQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_AX = CLBLM_L_X70Y124_SLICE_X104Y124_CO6;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C2 = CLBLM_L_X72Y114_SLICE_X109Y114_CO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D1 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D2 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D3 = 1'b1;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D4 = 1'b1;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C3 = CLBLM_L_X72Y118_SLICE_X108Y118_DO6;
  assign CLBLL_R_X75Y123_SLICE_X115Y123_D6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_BX = CLBLM_L_X70Y124_SLICE_X104Y124_AO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C1 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C2 = CLBLM_L_X70Y124_SLICE_X104Y124_AQ;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C4 = CLBLL_R_X73Y119_SLICE_X111Y119_CO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C3 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C5 = CLBLM_L_X70Y124_SLICE_X104Y124_BQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_C6 = RIOB33_X105Y161_IOB_X1Y161_I;
  assign CLBLM_L_X70Y119_SLICE_X104Y119_C5 = CLBLL_R_X73Y121_SLICE_X110Y121_CO6;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D1 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D2 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D3 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D4 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D5 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y87_ILOGIC_X1Y88_D = RIOB33_X105Y87_IOB_X1Y88_I;
  assign RIOI3_TBYTETERM_X105Y87_ILOGIC_X1Y87_D = RIOB33_X105Y87_IOB_X1Y87_I;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A1 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A2 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A3 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A4 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A5 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_A6 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B1 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B2 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B3 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B4 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B5 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_B6 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C1 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C2 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C3 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C4 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C5 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_C6 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D1 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D2 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D3 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D4 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D5 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X155Y131_D6 = 1'b1;
  assign LIOI3_X0Y159_ILOGIC_X0Y159_D = LIOB33_X0Y159_IOB_X0Y159_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A2 = RIOB33_X105Y187_IOB_X1Y187_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A3 = RIOB33_SING_X105Y199_IOB_X1Y199_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A5 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_A6 = RIOB33_SING_X105Y99_IOB_X1Y99_I;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B1 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B2 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B3 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B4 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B5 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_B6 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C1 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C2 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C3 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C4 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C5 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_C6 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D1 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D2 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D3 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D4 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D5 = 1'b1;
  assign CLBLM_L_X98Y131_SLICE_X154Y131_D6 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A3 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A4 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A5 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_A6 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B1 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B2 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B4 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B5 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C1 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C4 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C5 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_C6 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y157_D = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D1 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D3 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D5 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X75Y124_SLICE_X114Y124_D6 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A1 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A2 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A4 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A5 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_A6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B1 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B2 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B4 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B5 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_B6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C1 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C2 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C3 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C4 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_A1 = CLBLM_L_X72Y114_SLICE_X109Y114_CO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_A2 = CLBLL_R_X73Y121_SLICE_X110Y121_CO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_A3 = CLBLM_L_X72Y118_SLICE_X108Y118_DO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_A4 = CLBLL_R_X73Y119_SLICE_X111Y119_CO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_A5 = CLBLM_L_X72Y118_SLICE_X108Y118_CO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_A6 = CLBLM_L_X70Y117_SLICE_X105Y117_AO6;
  assign CLBLM_L_X72Y131_SLICE_X109Y131_C5 = 1'b1;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A1 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A3 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A4 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_B3 = CLBLM_L_X72Y118_SLICE_X108Y118_DO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_B4 = CLBLM_L_X72Y118_SLICE_X108Y118_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_B1 = CLBLM_L_X72Y114_SLICE_X109Y114_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_B2 = CLBLL_R_X73Y121_SLICE_X110Y121_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B1 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_C1 = CLBLL_R_X73Y119_SLICE_X111Y119_CO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_C2 = CLBLM_L_X70Y117_SLICE_X105Y117_AO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_C3 = CLBLL_R_X73Y121_SLICE_X110Y121_CO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_C4 = CLBLM_L_X72Y114_SLICE_X109Y114_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B2 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B3 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B4 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C1 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C2 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C5 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_C6 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_D1 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_D2 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_D3 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_D6 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_D4 = 1'b1;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_D5 = 1'b1;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D1 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D2 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D5 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X75Y124_SLICE_X115Y124_D6 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_A1 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_A2 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_A3 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_A4 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_A5 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_A6 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_B1 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_B2 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_B3 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_B4 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_B5 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_B6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D1 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D2 = CLBLM_L_X72Y128_SLICE_X109Y128_CO6;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D3 = CLBLM_L_X74Y128_SLICE_X112Y128_CO6;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_C1 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_C2 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_C3 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_C4 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_C5 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_C6 = 1'b1;
  assign CLBLM_L_X72Y131_SLICE_X108Y131_D6 = CLBLL_R_X75Y127_SLICE_X114Y127_CO6;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_D1 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_D2 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_D3 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_D4 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_D5 = 1'b1;
  assign CLBLM_L_X68Y119_SLICE_X102Y119_D6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A2 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A3 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A4 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A5 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_A6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B2 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B3 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B4 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B5 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_B6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C2 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C3 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C4 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C5 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_C6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D2 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D3 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D4 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D5 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X155Y132_D6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A4 = RIOB33_X105Y197_IOB_X1Y198_I;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A5 = RIOB33_X105Y185_IOB_X1Y186_I;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_A6 = RIOB33_X105Y97_IOB_X1Y98_I;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B2 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B3 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B4 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B5 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_B6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C2 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C3 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C4 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C5 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_C6 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D1 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D2 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D3 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D4 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D5 = 1'b1;
  assign CLBLM_L_X98Y132_SLICE_X154Y132_D6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_L_X70Y123_SLICE_X105Y123_DO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_A2 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_A3 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_A4 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_A5 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_B1 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_B2 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_B3 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_B5 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_C1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_C2 = CLBLL_R_X75Y125_SLICE_X115Y125_F7AMUX_O;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_C3 = CLBLM_L_X76Y125_SLICE_X116Y125_F8MUX_O;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_C4 = CLBLL_R_X75Y125_SLICE_X114Y125_F7AMUX_O;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_C5 = CLBLM_L_X70Y121_SLICE_X105Y121_CO6;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_C6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_D1 = 1'b1;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_D2 = 1'b1;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_D3 = 1'b1;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_D4 = 1'b1;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_D5 = 1'b1;
  assign CLBLL_R_X75Y125_SLICE_X114Y125_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLM_L_X70Y121_SLICE_X104Y121_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLM_L_X56Y116_SLICE_X84Y116_CO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_A2 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_A3 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_A4 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_A5 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_B1 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_B2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_B4 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_B6 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_C1 = CLBLL_R_X75Y126_SLICE_X115Y126_F7BMUX_O;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_C2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_C3 = CLBLL_R_X75Y126_SLICE_X115Y126_F7AMUX_O;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_C4 = CLBLM_L_X76Y125_SLICE_X117Y125_F8MUX_O;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_C5 = CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_A4 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_A5 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_D1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_D2 = CLBLM_L_X76Y124_SLICE_X116Y124_F7AMUX_O;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_D3 = CLBLL_R_X77Y125_SLICE_X118Y125_F8MUX_O;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_D4 = CLBLM_L_X70Y122_SLICE_X104Y122_CO6;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_D5 = CLBLM_L_X76Y124_SLICE_X116Y124_F7BMUX_O;
  assign CLBLL_R_X75Y125_SLICE_X115Y125_D6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_A1 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_A2 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_A3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_A4 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_A5 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_B2 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_B3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_B4 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_B5 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_B6 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_C1 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_C2 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_C4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_C6 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_D1 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_D2 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_D4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_D5 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X73Y114_SLICE_X110Y114_D6 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign LIOI3_X0Y183_ILOGIC_X0Y184_D = LIOB33_X0Y183_IOB_X0Y184_I;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D6 = CLBLM_L_X74Y117_SLICE_X113Y117_CO6;
  assign LIOI3_X0Y183_ILOGIC_X0Y183_D = LIOB33_X0Y183_IOB_X0Y183_I;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_A1 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_A2 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_A3 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_A4 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_A5 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_A6 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_B1 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_B2 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_B3 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_B4 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_B5 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_B6 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_C6 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_C1 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_C2 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_C3 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_C4 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_C5 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_C6 = 1'b1;
  assign RIOI3_X105Y167_ILOGIC_X1Y167_D = RIOB33_X105Y167_IOB_X1Y167_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_D1 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_D2 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_D3 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_D4 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_D5 = 1'b1;
  assign CLBLL_R_X73Y114_SLICE_X111Y114_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_A1 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_A2 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_A3 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_A4 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_A5 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_A6 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_B1 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_B2 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_B3 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_B4 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_B5 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_B6 = 1'b1;
  assign LIOB33_X0Y85_IOB_X0Y86_O = CLBLM_L_X70Y119_SLICE_X104Y119_AO6;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_C1 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_C2 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_C3 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_C4 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_C5 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_C6 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_D1 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_D2 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_D3 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_D4 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_D5 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X114Y126_D6 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_A1 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_A2 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_A3 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_A4 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_A5 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_A6 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_B1 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_B2 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_B3 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_B4 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_B5 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_B6 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_A2 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_A3 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D5 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_C1 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_C2 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_C3 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_C4 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_C5 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_C6 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_B2 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_B3 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_B4 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_B5 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_C1 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_C2 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_C3 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_D3 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_D4 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_D5 = 1'b1;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_D6 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y127_SLICE_X105Y127_D1 = 1'b1;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_D1 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_D2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_D4 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_D5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X75Y126_SLICE_X115Y126_D6 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_A1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_A2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_A3 = CLBLL_R_X73Y122_SLICE_X110Y122_DO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_A4 = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_A5 = CLBLM_L_X70Y128_SLICE_X104Y128_AO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_A6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_AX = CLBLM_L_X70Y127_SLICE_X104Y127_DO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_B1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_B3 = CLBLM_L_X70Y127_SLICE_X104Y127_AQ;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_B4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_B5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_B6 = CLBLM_L_X70Y127_SLICE_X104Y127_CO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_B2 = CLBLL_R_X71Y125_SLICE_X106Y125_BO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_A2 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_BX = CLBLM_L_X70Y127_SLICE_X104Y127_AO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_A3 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_C1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_C2 = CLBLM_L_X70Y127_SLICE_X104Y127_CQ;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_C3 = CLBLM_L_X70Y127_SLICE_X104Y127_AQ;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_C4 = RIOB33_X105Y183_IOB_X1Y184_I;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_C5 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_C6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_A5 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_A6 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_B2 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_B3 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_CX = CLBLM_L_X70Y127_SLICE_X104Y127_BO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_B4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_D1 = RIOB33_X105Y185_IOB_X1Y185_I;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_D2 = CLBLM_L_X70Y127_SLICE_X104Y127_CQ;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_D3 = CLBLM_L_X70Y127_SLICE_X104Y127_AQ;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_D4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_D5 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y127_SLICE_X104Y127_D6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_C2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_C3 = CLBLL_R_X73Y115_SLICE_X111Y115_F8MUX_O;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_C4 = CLBLL_R_X73Y115_SLICE_X110Y115_F7AMUX_O;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_C5 = CLBLM_L_X72Y115_SLICE_X109Y115_F7AMUX_O;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_C6 = CLBLL_R_X71Y119_SLICE_X106Y119_AO6;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_D1 = 1'b1;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_D2 = 1'b1;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_D3 = 1'b1;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_D4 = 1'b1;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_D5 = 1'b1;
  assign CLBLL_R_X73Y115_SLICE_X110Y115_D6 = 1'b1;
  assign LIOI3_X0Y173_ILOGIC_X0Y174_D = LIOB33_X0Y173_IOB_X0Y174_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y173_ILOGIC_X0Y173_D = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_A2 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_A2 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_A3 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_A4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_A6 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_B2 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_B3 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_B4 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_B5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_B6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_C1 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_C2 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_C3 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_C4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_C5 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_C6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_D1 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_D2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_D3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_D4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_D5 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X73Y115_SLICE_X111Y115_D6 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLM_R_X59Y117_SLICE_X88Y117_AO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_B1 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_B3 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_B4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_B5 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_B6 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign LIOB33_X0Y87_IOB_X0Y88_O = CLBLM_L_X70Y128_SLICE_X105Y128_AO6;
  assign LIOB33_X0Y87_IOB_X0Y87_O = CLBLL_R_X71Y119_SLICE_X106Y119_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A1 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A2 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_A6 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_C3 = CLBLL_R_X75Y115_SLICE_X115Y115_F8MUX_O;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B1 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B2 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B4 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B5 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_A6 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C1 = CLBLM_L_X70Y122_SLICE_X104Y122_CO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C3 = CLBLL_R_X75Y127_SLICE_X115Y127_F8MUX_O;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C4 = CLBLL_R_X75Y127_SLICE_X114Y127_F7AMUX_O;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C5 = CLBLM_L_X74Y127_SLICE_X113Y127_F7AMUX_O;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y116_SLICE_X114Y116_C6 = CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D1 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D2 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D3 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D4 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D5 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X114Y127_D6 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A1 = CLBLM_L_X70Y128_SLICE_X105Y128_AQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A2 = CLBLL_R_X71Y127_SLICE_X106Y127_AO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A3 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A4 = CLBLM_L_X70Y128_SLICE_X105Y128_BO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A1 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A2 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A4 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A5 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_A6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_A6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_AX = CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B2 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B4 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B5 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_B6 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B2 = CLBLM_L_X70Y128_SLICE_X105Y128_BQ;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B3 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C1 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C2 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C3 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_C6 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C6 = RIOB33_X105Y153_IOB_X1Y153_I;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_C4 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D1 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D2 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D3 = 1'b1;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D1 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D2 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D4 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D5 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X75Y127_SLICE_X115Y127_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D4 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A2 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A3 = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A4 = CLBLM_L_X70Y127_SLICE_X104Y127_BQ;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_A6 = RIOB33_X105Y179_IOB_X1Y180_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_L_X70Y127_SLICE_X104Y127_BO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_AX = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B1 = RIOB33_X105Y181_IOB_X1Y181_I;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_A1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_A2 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_A3 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_A5 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_A6 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B2 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B3 = CLBLM_L_X70Y128_SLICE_X104Y128_AQ;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_B4 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_B1 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_B2 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_B3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_B4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_B5 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C1 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_C2 = 1'b1;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_C1 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_C2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_C3 = CLBLL_R_X73Y116_SLICE_X111Y116_F8MUX_O;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_C4 = CLBLL_R_X73Y116_SLICE_X110Y116_F7AMUX_O;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_C5 = CLBLM_L_X72Y116_SLICE_X109Y116_F7BMUX_O;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D1 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D2 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D3 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D4 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D5 = 1'b1;
  assign CLBLM_L_X70Y128_SLICE_X104Y128_D6 = 1'b1;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_D1 = 1'b1;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_D2 = 1'b1;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_D3 = 1'b1;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_D4 = 1'b1;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_D5 = 1'b1;
  assign CLBLL_R_X73Y116_SLICE_X110Y116_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_L_X70Y121_SLICE_X104Y121_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_A1 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_A3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_A4 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_A5 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_A6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_B1 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_B3 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_B4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_B5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_B6 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_C1 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_C2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_C3 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_C4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_C5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_C6 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_D1 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_D2 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_D4 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_D5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y116_SLICE_X111Y116_D6 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_A3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOB33_X0Y89_IOB_X0Y90_O = CLBLL_R_X71Y128_SLICE_X106Y128_AO6;
  assign LIOB33_X0Y89_IOB_X0Y89_O = CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  assign LIOI3_X0Y185_ILOGIC_X0Y186_D = LIOB33_X0Y185_IOB_X0Y186_I;
  assign LIOI3_X0Y185_ILOGIC_X0Y185_D = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A1 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A2 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A5 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_A6 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B2 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B4 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_B6 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C2 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C3 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C4 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C5 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_C6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign RIOI3_X105Y171_ILOGIC_X1Y172_D = RIOB33_X105Y171_IOB_X1Y172_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y171_ILOGIC_X1Y171_D = RIOB33_X105Y171_IOB_X1Y171_I;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D3 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D4 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D5 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X75Y128_SLICE_X114Y128_D6 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A1 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A2 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_A6 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A1 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A2 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_A3 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B1 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B3 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B5 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_B6 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_B1 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C2 = CLBLM_L_X76Y127_SLICE_X116Y127_F7AMUX_O;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C3 = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C4 = CLBLL_R_X75Y128_SLICE_X115Y128_F7AMUX_O;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C5 = CLBLM_L_X76Y128_SLICE_X116Y128_F8MUX_O;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C1 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C2 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C3 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C4 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C5 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_C6 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D1 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D2 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D3 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D4 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D5 = 1'b1;
  assign CLBLL_R_X75Y128_SLICE_X115Y128_D6 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D1 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D2 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D3 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D4 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D5 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X105Y129_D6 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A1 = CLBLM_L_X70Y129_SLICE_X104Y129_BO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A3 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A4 = CLBLL_R_X71Y129_SLICE_X106Y129_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A5 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_A6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_AX = CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B2 = CLBLM_L_X70Y129_SLICE_X104Y129_BQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B3 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B5 = RIOB33_X105Y157_IOB_X1Y158_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_B6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_BX = CLBLM_L_X70Y129_SLICE_X104Y129_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C1 = CLBLM_L_X70Y129_SLICE_X104Y129_BQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C2 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C3 = CLBLM_L_X70Y129_SLICE_X104Y129_AQ;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C4 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C5 = RIOB33_X105Y159_IOB_X1Y159_I;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_C6 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D1 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D2 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D3 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D4 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D5 = 1'b1;
  assign CLBLM_L_X70Y129_SLICE_X104Y129_D6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_B6 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C4 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C5 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X113Y120_C6 = 1'b1;
  assign LIOB33_X0Y91_IOB_X0Y92_O = CLBLL_R_X71Y131_SLICE_X107Y131_BO6;
  assign LIOB33_X0Y91_IOB_X0Y91_O = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_C2 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_C3 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_C4 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_C5 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B5 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_B6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A2 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A3 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A4 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_A6 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B2 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B3 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B5 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C2 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C4 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_C6 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D1 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D2 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D4 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y118_SLICE_X110Y118_D6 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C5 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_L_X74Y120_SLICE_X112Y120_C6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A2 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A5 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_A6 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B1 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B2 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B3 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B5 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C1 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C2 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C3 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C4 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C5 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_C6 = 1'b1;
  assign LIOB33_X0Y93_IOB_X0Y94_O = CLBLM_L_X70Y129_SLICE_X104Y129_AO6;
  assign LIOB33_X0Y93_IOB_X0Y93_O = CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D1 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D2 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D3 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D4 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D5 = 1'b1;
  assign CLBLL_R_X73Y118_SLICE_X111Y118_D6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_B6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_L_X70Y127_SLICE_X104Y127_DO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C1 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B2 = 1'b1;
  assign CLBLM_L_X74Y129_SLICE_X112Y129_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C2 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_B3 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C3 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X117Y127_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C1 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_C2 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D1 = 1'b1;
  assign CLBLL_R_X77Y129_SLICE_X119Y129_D4 = 1'b1;
  assign LIOI3_X0Y189_ILOGIC_X0Y190_D = LIOB33_X0Y189_IOB_X0Y190_I;
  assign LIOI3_X0Y189_ILOGIC_X0Y189_D = LIOB33_X0Y189_IOB_X0Y189_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A1 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A3 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A5 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_A6 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B1 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B3 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B4 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C2 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C4 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C5 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_C6 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y173_ILOGIC_X1Y174_D = RIOB33_X105Y173_IOB_X1Y174_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y173_ILOGIC_X1Y173_D = RIOB33_X105Y173_IOB_X1Y173_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D1 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D4 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D5 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X73Y119_SLICE_X110Y119_D6 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B2 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y51_ILOGIC_X1Y52_D = RIOB33_X105Y51_IOB_X1Y52_I;
  assign RIOI3_X105Y51_ILOGIC_X1Y51_D = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_B6 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y164_D = RIOB33_X105Y163_IOB_X1Y164_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A3 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A4 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_A6 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign LIOB33_X0Y95_IOB_X0Y95_O = CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  assign LIOB33_X0Y95_IOB_X0Y96_O = CLBLM_L_X70Y124_SLICE_X104Y124_AO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign RIOI3_TBYTETERM_X105Y163_ILOGIC_X1Y163_D = RIOB33_X105Y163_IOB_X1Y163_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B2 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B3 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B5 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_B6 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C1 = CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C4 = CLBLL_R_X73Y119_SLICE_X111Y119_F7AMUX_O;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C5 = CLBLL_R_X73Y118_SLICE_X111Y118_F7AMUX_O;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_C6 = CLBLM_L_X74Y119_SLICE_X112Y119_F8MUX_O;
  assign RIOI3_TBYTESRC_X105Y57_ILOGIC_X1Y57_D = RIOB33_X105Y57_IOB_X1Y57_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C1 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C2 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D3 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D4 = 1'b1;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X73Y119_SLICE_X111Y119_D6 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C5 = 1'b1;
  assign CLBLM_L_X76Y127_SLICE_X116Y127_C6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_A1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_A3 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_A4 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_A6 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_B1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_B2 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_B3 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_B5 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_C2 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_C3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_C4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_C5 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_C6 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_D1 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_D2 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_D3 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_D4 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_D5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y120_SLICE_X110Y120_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOB33_X0Y97_IOB_X0Y98_O = CLBLL_R_X71Y131_SLICE_X106Y131_AO6;
  assign LIOB33_X0Y97_IOB_X0Y97_O = CLBLM_L_X70Y124_SLICE_X104Y124_CO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_A1 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_A2 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_A3 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_A5 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_A6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_B1 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_B3 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_B4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_B5 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_C1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_C2 = CLBLL_R_X73Y120_SLICE_X110Y120_F7AMUX_O;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_C3 = CLBLL_R_X75Y120_SLICE_X114Y120_F8MUX_O;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_C4 = CLBLL_R_X73Y120_SLICE_X110Y120_F7BMUX_O;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_C5 = CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_C6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_D3 = CLBLL_R_X73Y120_SLICE_X111Y120_DO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_D4 = CLBLM_L_X72Y120_SLICE_X108Y120_DO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_D1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_D2 = CLBLL_R_X73Y121_SLICE_X111Y121_F7AMUX_O;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_D3 = CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_D4 = CLBLL_R_X73Y120_SLICE_X111Y120_F7AMUX_O;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_D5 = CLBLM_L_X74Y120_SLICE_X112Y120_F8MUX_O;
  assign CLBLL_R_X73Y120_SLICE_X111Y120_D6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_A6 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign RIOI3_X105Y165_ILOGIC_X1Y166_D = RIOB33_X105Y165_IOB_X1Y166_I;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y117_SLICE_X114Y117_B6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign RIOI3_X105Y165_ILOGIC_X1Y165_D = RIOB33_X105Y165_IOB_X1Y165_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_D4 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_D5 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A2 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A3 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A4 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_A6 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C2 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B1 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B3 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B5 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_B6 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C3 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C1 = CLBLM_L_X70Y129_SLICE_X104Y129_CO6;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C2 = CLBLL_R_X73Y121_SLICE_X111Y121_F7BMUX_O;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C3 = CLBLM_L_X74Y121_SLICE_X112Y121_F8MUX_O;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C4 = CLBLL_R_X73Y121_SLICE_X110Y121_F7AMUX_O;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y126_SLICE_X109Y126_C5 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_A4 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLM_R_X59Y117_SLICE_X88Y117_AO6;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D1 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D2 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D3 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D4 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D5 = 1'b1;
  assign CLBLL_R_X73Y121_SLICE_X110Y121_D6 = 1'b1;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_A6 = CLBLL_R_X71Y116_SLICE_X107Y116_DO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_AX = CLBLM_L_X70Y121_SLICE_X105Y121_CO6;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D1 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A2 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_A6 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_C3 = CLBLL_R_X75Y118_SLICE_X115Y118_F8MUX_O;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B2 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B4 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B5 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_B6 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C1 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C2 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C3 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_C6 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D2 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D3 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D4 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y121_SLICE_X111Y121_D6 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign LIOI3_X0Y191_ILOGIC_X0Y192_D = LIOB33_X0Y191_IOB_X0Y192_I;
  assign LIOI3_X0Y191_ILOGIC_X0Y191_D = LIOB33_X0Y191_IOB_X0Y191_I;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_C3 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign RIOI3_X105Y175_ILOGIC_X1Y176_D = RIOB33_X105Y175_IOB_X1Y176_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign RIOI3_X105Y175_ILOGIC_X1Y175_D = RIOB33_X105Y175_IOB_X1Y175_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y53_ILOGIC_X1Y54_D = RIOB33_X105Y53_IOB_X1Y54_I;
  assign RIOI3_X105Y53_ILOGIC_X1Y53_D = RIOB33_X105Y53_IOB_X1Y53_I;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_D2 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y188_D = RIOB33_X105Y187_IOB_X1Y188_I;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D6 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign RIOI3_TBYTETERM_X105Y187_ILOGIC_X1Y187_D = RIOB33_X105Y187_IOB_X1Y187_I;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_D4 = 1'b1;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_D5 = 1'b1;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign RIOI3_TBYTESRC_X105Y69_ILOGIC_X1Y70_D = RIOB33_X105Y69_IOB_X1Y70_I;
  assign CLBLM_L_X70Y121_SLICE_X105Y121_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y69_ILOGIC_X1Y69_D = RIOB33_X105Y69_IOB_X1Y69_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_A2 = CLBLM_L_X70Y123_SLICE_X104Y123_AO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_A3 = CLBLM_L_X70Y121_SLICE_X104Y121_AQ;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_A4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_AX = CLBLM_L_X70Y123_SLICE_X104Y123_BO6;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_B1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A1 = CLBLL_R_X73Y123_SLICE_X110Y123_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A2 = CLBLL_R_X73Y123_SLICE_X110Y123_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A3 = CLBLM_L_X74Y125_SLICE_X112Y125_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A4 = CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A5 = CLBLM_L_X74Y123_SLICE_X112Y123_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_A6 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_B2 = CLBLM_L_X70Y121_SLICE_X104Y121_BQ;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_B3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B1 = CLBLL_R_X73Y123_SLICE_X110Y123_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B2 = CLBLL_R_X73Y123_SLICE_X110Y123_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B3 = CLBLM_L_X74Y123_SLICE_X112Y123_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B4 = CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B5 = CLBLM_L_X74Y125_SLICE_X112Y125_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_B6 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_B4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_B5 = CLBLM_L_X70Y121_SLICE_X104Y121_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C1 = CLBLM_L_X74Y125_SLICE_X112Y125_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C2 = CLBLM_L_X74Y123_SLICE_X112Y123_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C3 = CLBLL_R_X73Y123_SLICE_X110Y123_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C4 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C5 = CLBLL_R_X73Y123_SLICE_X110Y123_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_C6 = CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_B6 = CLBLM_L_X72Y120_SLICE_X108Y120_CO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D2 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D3 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D1 = CLBLM_L_X74Y125_SLICE_X112Y125_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D2 = CLBLL_R_X75Y123_SLICE_X114Y123_AO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D3 = CLBLL_R_X73Y123_SLICE_X110Y123_DO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D4 = CLBLM_L_X74Y123_SLICE_X112Y123_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D5 = CLBLL_R_X73Y123_SLICE_X110Y123_CO6;
  assign CLBLL_R_X73Y122_SLICE_X110Y122_D6 = CLBLM_L_X72Y122_SLICE_X108Y122_AO6;
  assign CLBLM_L_X72Y126_SLICE_X108Y126_D4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_BX = CLBLM_L_X70Y121_SLICE_X104Y121_DO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_C2 = CLBLM_L_X70Y121_SLICE_X104Y121_CQ;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_C3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A1 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A2 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A3 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A4 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A5 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_A6 = 1'b1;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_C5 = RIOB33_X105Y177_IOB_X1Y178_I;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_C6 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B1 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B2 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B3 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B4 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B5 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_B6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B5 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C1 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C2 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C3 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C4 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C5 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_C6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_B6 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X70Y121_SLICE_X104Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D1 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D2 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D3 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D4 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D5 = 1'b1;
  assign CLBLL_R_X73Y122_SLICE_X111Y122_D6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_C6 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A3 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A4 = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A6 = CLBLL_R_X71Y118_SLICE_X106Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_AX = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B2 = CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B3 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B5 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D5 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X74Y121_SLICE_X113Y121_D6 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_BX = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C1 = CLBLL_L_X2Y118_SLICE_X0Y118_BQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C2 = CLBLL_L_X2Y118_SLICE_X0Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C3 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C6 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_L_X70Y119_SLICE_X105Y119_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D6 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_A6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A2 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y124_SLICE_X116Y124_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A4 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A5 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_B1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_A6 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_CE = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D6 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A1 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A3 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_A6 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B3 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B4 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B5 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_B6 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B2 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B3 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C2 = CLBLM_L_X74Y123_SLICE_X112Y123_F7AMUX_O;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C3 = CLBLL_R_X73Y123_SLICE_X111Y123_F8MUX_O;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C4 = CLBLL_R_X73Y123_SLICE_X110Y123_F7AMUX_O;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_C6 = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B4 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_C3 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_B6 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_C4 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D2 = CLBLL_R_X73Y124_SLICE_X111Y124_F7AMUX_O;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D3 = CLBLM_L_X74Y124_SLICE_X112Y124_F8MUX_O;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D4 = CLBLL_R_X73Y124_SLICE_X111Y124_F7BMUX_O;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y123_SLICE_X110Y123_D6 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_C5 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_C6 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C1 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C3 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A2 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A3 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A4 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A5 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B1 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B2 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B3 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_B6 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_C6 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C2 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C3 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C4 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C5 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_C6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D1 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D2 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D4 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D5 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X73Y123_SLICE_X111Y123_D6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D5 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLM_L_X74Y121_SLICE_X112Y121_D6 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_B3 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = CLBLM_L_X68Y119_SLICE_X103Y119_BO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_AX = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = CLBLL_L_X2Y119_SLICE_X0Y119_BQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C1 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_C2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_BX = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = CLBLL_L_X2Y119_SLICE_X0Y119_AQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = CLBLL_L_X2Y119_SLICE_X0Y119_BQ;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_B4 = RIOB33_X105Y75_IOB_X1Y75_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_B5 = RIOB33_X105Y191_IOB_X1Y191_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_B6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y196_D = LIOB33_X0Y195_IOB_X0Y196_I;
  assign LIOI3_X0Y195_ILOGIC_X0Y195_D = LIOB33_X0Y195_IOB_X0Y195_I;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLM_L_X70Y121_SLICE_X104Y121_AO6;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLM_L_X56Y116_SLICE_X84Y116_CO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D1 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_C1 = 1'b1;
  assign RIOI3_X105Y177_ILOGIC_X1Y178_D = RIOB33_X105Y177_IOB_X1Y178_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = CLBLM_L_X68Y119_SLICE_X103Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_AX = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = CLBLL_L_X2Y119_SLICE_X1Y119_BQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D5 = 1'b1;
  assign CLBLL_R_X77Y130_SLICE_X119Y130_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_BX = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLM_L_X76Y128_SLICE_X117Y128_D6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = CLBLL_L_X2Y119_SLICE_X1Y119_BQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_C6 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y55_ILOGIC_X1Y56_D = RIOB33_X105Y55_IOB_X1Y56_I;
  assign LIOI3_TBYTESRC_X0Y157_ILOGIC_X0Y158_D = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = 1'b1;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A1 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A2 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A5 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_A6 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B1 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B4 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B5 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_B6 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C1 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C2 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C5 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_C6 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A2 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign RIOI3_TBYTESRC_X105Y81_ILOGIC_X1Y82_D = RIOB33_X105Y81_IOB_X1Y82_I;
  assign RIOI3_TBYTESRC_X105Y81_ILOGIC_X1Y81_D = RIOB33_X105Y81_IOB_X1Y81_I;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D1 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D2 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X73Y124_SLICE_X110Y124_D6 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A4 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A5 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_A6 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_D4 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_D5 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_D6 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A1 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A2 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A4 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A5 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B1 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B2 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B4 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B2 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B3 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C1 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C2 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C3 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C5 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_C6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B5 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_B6 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D1 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D2 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X73Y124_SLICE_X111Y124_D6 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C1 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C2 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C4 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_C6 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_A1 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_A3 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_A4 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_A5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_A6 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_B1 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_B3 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_B4 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_B5 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_B6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y182_D = LIOB33_X0Y181_IOB_X0Y182_I;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_C1 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_C2 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_C3 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_C4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_C6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = CLBLL_R_X71Y119_SLICE_X106Y119_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = CLBLL_L_X2Y120_SLICE_X0Y120_AQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_D1 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_AX = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_D2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = CLBLL_L_X2Y120_SLICE_X0Y120_BQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = CLBLL_L_X2Y120_SLICE_X0Y120_AQ;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_D4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_BX = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_R_X71Y116_SLICE_X106Y116_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = CLBLL_L_X2Y120_SLICE_X0Y120_BQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = CLBLL_L_X2Y120_SLICE_X0Y120_AQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D3 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLM_L_X70Y123_SLICE_X104Y123_BO6;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_L_X70Y123_SLICE_X105Y123_AO6;
  assign CLBLM_L_X76Y128_SLICE_X116Y128_D5 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_A1 = CLBLM_L_X72Y116_SLICE_X108Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_A2 = CLBLM_L_X74Y116_SLICE_X113Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_A3 = CLBLM_L_X72Y119_SLICE_X108Y119_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_A4 = CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_A5 = CLBLL_R_X73Y115_SLICE_X110Y115_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_A6 = CLBLL_R_X75Y116_SLICE_X114Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_B1 = CLBLM_L_X72Y116_SLICE_X108Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_B2 = CLBLM_L_X74Y116_SLICE_X113Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_B3 = CLBLM_L_X72Y119_SLICE_X108Y119_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_B4 = CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_B5 = CLBLL_R_X73Y115_SLICE_X110Y115_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_B6 = CLBLL_R_X75Y116_SLICE_X114Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_C1 = CLBLL_R_X73Y115_SLICE_X110Y115_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_C2 = CLBLM_L_X74Y116_SLICE_X113Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_C3 = CLBLM_L_X72Y116_SLICE_X108Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_C4 = CLBLM_L_X72Y119_SLICE_X108Y119_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_C5 = CLBLL_R_X75Y116_SLICE_X114Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_C6 = CLBLM_L_X72Y119_SLICE_X108Y119_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = 1'b1;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_D1 = CLBLL_R_X73Y115_SLICE_X110Y115_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_D5 = CLBLL_R_X75Y116_SLICE_X114Y116_CO6;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_D2 = CLBLM_L_X74Y116_SLICE_X113Y116_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = 1'b1;
  assign CLBLL_R_X71Y116_SLICE_X107Y116_D6 = CLBLM_L_X72Y116_SLICE_X108Y116_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = 1'b1;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A2 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A3 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A4 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_A6 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B1 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B2 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B3 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C2 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C3 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C5 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_C6 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D1 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D2 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D3 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D4 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y125_SLICE_X110Y125_D6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A1 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A3 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A4 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_A6 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B4 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B5 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_B6 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C1 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C3 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C4 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_C6 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign RIOI3_X105Y55_ILOGIC_X1Y55_D = RIOB33_X105Y55_IOB_X1Y55_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D1 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D2 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D4 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D5 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X73Y125_SLICE_X111Y125_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A1 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A2 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A5 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_A6 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B1 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B2 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B5 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_B6 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C3 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C5 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_C6 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_L_X72Y131_SLICE_X108Y131_AO6;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLM_L_X70Y123_SLICE_X105Y123_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A3 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A4 = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A5 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A6 = CLBLM_L_X68Y119_SLICE_X103Y119_AO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D3 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D4 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D6 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y117_SLICE_X106Y117_D2 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B4 = CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B5 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B6 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C2 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C4 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C5 = CLBLL_L_X2Y123_SLICE_X0Y123_DQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C6 = CLBLL_L_X2Y123_SLICE_X0Y123_BQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_C5 = CLBLL_R_X75Y119_SLICE_X114Y119_F7AMUX_O;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_C6 = CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D1 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D2 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D3 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D5 = CLBLL_L_X2Y123_SLICE_X0Y123_DQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D6 = CLBLL_L_X2Y123_SLICE_X0Y123_BQ;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A2 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_A6 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B2 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_B6 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A4 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C2 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_C6 = 1'b1;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_A5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A6 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D3 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D4 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D1 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D5 = 1'b1;
  assign CLBLL_R_X71Y117_SLICE_X107Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_ILOGIC_X0Y181_D = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLL_R_X75Y118_SLICE_X114Y118_D6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D6 = 1'b1;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A2 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A3 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A4 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_A6 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B1 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B2 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B4 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C2 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C3 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C4 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_C6 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X70Y128_SLICE_X105Y128_D6 = 1'b1;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D3 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D4 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D5 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X73Y126_SLICE_X110Y126_D6 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_C3 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign LIOI3_X0Y197_ILOGIC_X0Y198_D = LIOB33_X0Y197_IOB_X0Y198_I;
  assign LIOI3_X0Y197_ILOGIC_X0Y197_D = LIOB33_X0Y197_IOB_X0Y197_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A1 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A5 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_A6 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B2 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B4 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_B6 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y179_ILOGIC_X1Y180_D = RIOB33_X105Y179_IOB_X1Y180_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C1 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C2 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C5 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_C6 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign RIOI3_X105Y179_ILOGIC_X1Y179_D = RIOB33_X105Y179_IOB_X1Y179_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D2 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D3 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D4 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y126_SLICE_X111Y126_D6 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y59_ILOGIC_X1Y60_D = RIOB33_X105Y59_IOB_X1Y60_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y170_D = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D2 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign RIOI3_X105Y59_ILOGIC_X1Y59_D = RIOB33_X105Y59_IOB_X1Y59_I;
  assign LIOI3_TBYTESRC_X0Y169_ILOGIC_X0Y169_D = LIOB33_X0Y169_IOB_X0Y169_I;
  assign CLBLM_L_X72Y127_SLICE_X109Y127_D3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign RIOI3_SING_X105Y150_ILOGIC_X1Y150_D = RIOB33_SING_X105Y150_IOB_X1Y150_I;
  assign RIOI3_TBYTESRC_X105Y93_ILOGIC_X1Y94_D = RIOB33_X105Y93_IOB_X1Y94_I;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign RIOI3_TBYTESRC_X105Y93_ILOGIC_X1Y93_D = RIOB33_X105Y93_IOB_X1Y93_I;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_A3 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_A4 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y118_SLICE_X115Y118_A6 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_A1 = CLBLM_L_X74Y117_SLICE_X113Y117_DO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_A2 = CLBLL_R_X75Y118_SLICE_X114Y118_CO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_A3 = CLBLM_L_X74Y117_SLICE_X113Y117_CO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_A4 = CLBLL_R_X73Y116_SLICE_X110Y116_CO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_A5 = CLBLM_L_X72Y116_SLICE_X108Y116_DO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_A6 = CLBLL_R_X75Y120_SLICE_X115Y120_CO6;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLL_R_X71Y131_SLICE_X107Y131_AO6;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_L_X70Y122_SLICE_X104Y122_AO6;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_B1 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_B2 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_B3 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_B4 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_B5 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_B6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_C1 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_C2 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_C3 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_C4 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_C5 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_C6 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_D1 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_D2 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_D3 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_D4 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_D5 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X106Y118_D6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOB33_SING_X0Y99_IOB_X0Y99_O = CLBLL_R_X71Y131_SLICE_X106Y131_CO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_A1 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_A2 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_A4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_A5 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_A6 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_A1 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_A2 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_B1 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_B3 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_B4 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_B5 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_A6 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_B1 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_C2 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_C3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_C4 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_C5 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_C6 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_B2 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_B3 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_B4 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_B5 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_B6 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_C1 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_C2 = 1'b1;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_D2 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_D3 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_D4 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_D5 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X71Y118_SLICE_X107Y118_D6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_C6 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_D1 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_D2 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_D3 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_D4 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_D5 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_D6 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_A2 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_A3 = LIOB33_X0Y161_IOB_X0Y161_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_A4 = RIOB33_X105Y55_IOB_X1Y55_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_A5 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_A6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A1 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A2 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A3 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_A6 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_B3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_B4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_B5 = LIOB33_X0Y155_IOB_X0Y155_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B2 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B4 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_B6 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_C1 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_C2 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C2 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C4 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C5 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_C6 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_D1 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_D2 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_D3 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_D4 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_D5 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_D6 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D2 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D3 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D5 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y127_SLICE_X110Y127_D6 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_B3 = CLBLM_L_X70Y122_SLICE_X104Y122_AQ;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_B4 = RIOB33_X105Y171_IOB_X1Y172_I;
  assign CLBLM_L_X70Y122_SLICE_X104Y122_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLM_R_X59Y118_SLICE_X88Y118_AO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A1 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A4 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_A6 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B2 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B5 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_B6 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C1 = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C2 = CLBLM_L_X74Y127_SLICE_X112Y127_F7AMUX_O;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C3 = CLBLL_R_X73Y127_SLICE_X110Y127_F8MUX_O;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C4 = CLBLL_R_X73Y127_SLICE_X111Y127_F7AMUX_O;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D1 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D2 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D3 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D4 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D5 = 1'b1;
  assign CLBLL_R_X73Y127_SLICE_X111Y127_D6 = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X70Y121_SLICE_X105Y121_AO6;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_L_X70Y122_SLICE_X104Y122_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A1 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A2 = RIOB33_X105Y151_IOB_X1Y151_I;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A3 = CLBLL_R_X71Y119_SLICE_X106Y119_AQ;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A4 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A5 = CLBLM_L_X70Y119_SLICE_X104Y119_AQ;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_A6 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B1 = CLBLM_L_X72Y116_SLICE_X108Y116_DO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B2 = CLBLM_L_X74Y117_SLICE_X113Y117_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B3 = CLBLL_R_X73Y116_SLICE_X110Y116_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B4 = CLBLL_R_X75Y118_SLICE_X114Y118_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B5 = CLBLM_L_X74Y117_SLICE_X113Y117_DO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_B6 = CLBLL_R_X75Y120_SLICE_X115Y120_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C1 = CLBLM_L_X74Y117_SLICE_X113Y117_DO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C2 = CLBLL_R_X75Y120_SLICE_X115Y120_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C3 = CLBLL_R_X73Y116_SLICE_X110Y116_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C4 = CLBLL_R_X75Y118_SLICE_X114Y118_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C5 = CLBLM_L_X72Y116_SLICE_X108Y116_DO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_C6 = CLBLM_L_X74Y117_SLICE_X113Y117_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A3 = CLBLL_L_X2Y123_SLICE_X0Y123_AQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A4 = CLBLL_L_X2Y123_SLICE_X0Y123_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_A6 = CLBLL_R_X71Y120_SLICE_X107Y120_BO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D3 = CLBLL_R_X73Y116_SLICE_X110Y116_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D4 = CLBLL_R_X75Y118_SLICE_X114Y118_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D1 = CLBLM_L_X74Y117_SLICE_X113Y117_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_AX = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D5 = CLBLM_L_X72Y116_SLICE_X108Y116_DO6;
  assign CLBLL_R_X71Y119_SLICE_X106Y119_D2 = CLBLL_R_X75Y120_SLICE_X115Y120_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B3 = CLBLL_L_X2Y123_SLICE_X0Y123_AQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B4 = CLBLL_L_X2Y123_SLICE_X0Y123_CQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B5 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_B6 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_BX = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C1 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C2 = CLBLL_L_X2Y123_SLICE_X0Y123_CQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C3 = CLBLL_L_X2Y123_SLICE_X0Y123_AQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C5 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_C6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_CX = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D1 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D2 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D3 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D4 = CLBLL_L_X2Y124_SLICE_X0Y124_AQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D5 = CLBLL_L_X2Y124_SLICE_X0Y124_CQ;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_D6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A1 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A2 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X0Y123_DX = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A3 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A4 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_A6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B1 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B2 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B4 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B5 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_B6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C1 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C4 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C5 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_C6 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A1 = CLBLL_L_X2Y124_SLICE_X1Y124_DQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A2 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A3 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A4 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A5 = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_A6 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D1 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D2 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B2 = CLBLL_L_X2Y124_SLICE_X0Y124_AQ;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_B6 = CLBLL_L_X2Y124_SLICE_X0Y124_CQ;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D4 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLL_R_X71Y119_SLICE_X107Y119_D6 = CLBLM_L_X78Y121_SLICE_X120Y121_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_C6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D1 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D2 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D3 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D4 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D5 = 1'b1;
  assign CLBLL_L_X2Y123_SLICE_X1Y123_D6 = 1'b1;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A2 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A4 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A5 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_A6 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B2 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B4 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B5 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_B6 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C1 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C2 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C3 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C4 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_C6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y177_ILOGIC_X1Y177_D = RIOB33_X105Y177_IOB_X1Y177_I;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D2 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D4 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D5 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X73Y128_SLICE_X110Y128_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A3 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A4 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_A6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B1 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B2 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B3 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_B6 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C2 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C3 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C4 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C5 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_C6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D1 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D4 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D5 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X73Y128_SLICE_X111Y128_D6 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_L_X70Y119_SLICE_X105Y119_AO6;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_L_X70Y121_SLICE_X105Y121_CO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_A1 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_A3 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_A4 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_A5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B1 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B2 = 1'b1;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y201_ILOGIC_X0Y202_D = LIOB33_X0Y201_IOB_X0Y202_I;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_B1 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_B2 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_B3 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_B4 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_B5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_B3 = 1'b1;
  assign LIOI3_X0Y201_ILOGIC_X0Y201_D = LIOB33_X0Y201_IOB_X0Y201_I;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_C1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_C2 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_C3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_C4 = CLBLL_R_X77Y129_SLICE_X118Y129_BO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_C5 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_C6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A2 = CLBLL_L_X2Y124_SLICE_X0Y124_BQ;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A4 = CLBLL_L_X2Y124_SLICE_X0Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A5 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_A6 = CLBLL_R_X71Y126_SLICE_X106Y126_AO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_D4 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_D1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_D6 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_AX = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_D5 = CLBLM_L_X78Y124_SLICE_X120Y124_BO6;
  assign CLBLL_R_X71Y120_SLICE_X106Y120_D2 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B3 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B5 = CLBLL_L_X2Y124_SLICE_X0Y124_BQ;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_B6 = CLBLL_L_X2Y124_SLICE_X0Y124_DQ;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_BX = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C1 = CLBLL_L_X2Y124_SLICE_X0Y124_BQ;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C2 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C3 = CLBLL_L_X2Y124_SLICE_X0Y124_DQ;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C5 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_C6 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C1 = 1'b1;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C2 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_CX = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D1 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D2 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D3 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D4 = CLBLL_L_X2Y124_SLICE_X1Y124_CQ;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D5 = CLBLL_L_X2Y124_SLICE_X1Y124_BQ;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_D6 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_A1 = CLBLM_L_X70Y127_SLICE_X104Y127_DO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y124_SLICE_X0Y124_DX = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_A3 = CLBLL_R_X71Y119_SLICE_X107Y119_F7BMUX_O;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_A4 = CLBLL_R_X71Y120_SLICE_X106Y120_F7AMUX_O;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_A6 = CLBLM_L_X72Y120_SLICE_X109Y120_F8MUX_O;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C6 = 1'b1;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_B1 = CLBLL_R_X73Y120_SLICE_X111Y120_CO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_B2 = CLBLM_L_X74Y120_SLICE_X113Y120_AO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_B3 = CLBLM_L_X72Y120_SLICE_X108Y120_DO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_B4 = CLBLL_R_X73Y120_SLICE_X111Y120_DO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_B5 = CLBLL_R_X71Y120_SLICE_X107Y120_AO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_B6 = CLBLL_R_X71Y122_SLICE_X106Y122_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A2 = 1'b1;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_C1 = CLBLL_R_X71Y120_SLICE_X107Y120_AO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_C2 = CLBLM_L_X74Y120_SLICE_X113Y120_AO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_C3 = CLBLM_L_X72Y120_SLICE_X108Y120_DO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_C4 = CLBLL_R_X71Y122_SLICE_X106Y122_AO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_C5 = CLBLL_R_X73Y120_SLICE_X111Y120_CO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_C6 = CLBLL_R_X73Y120_SLICE_X111Y120_DO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A3 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A4 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A5 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_A6 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A1 = CLBLL_R_X71Y125_SLICE_X106Y125_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A3 = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A4 = CLBLL_L_X2Y124_SLICE_X1Y124_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_A6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_D1 = CLBLL_R_X71Y120_SLICE_X107Y120_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_AX = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_D5 = CLBLL_R_X73Y120_SLICE_X111Y120_CO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_D2 = CLBLL_R_X71Y122_SLICE_X106Y122_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B3 = CLBLL_L_X2Y124_SLICE_X1Y124_AQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B5 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_B6 = CLBLL_L_X2Y124_SLICE_X1Y124_DQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_BX = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLL_R_X71Y120_SLICE_X107Y120_D6 = CLBLM_L_X74Y120_SLICE_X113Y120_AO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C2 = CLBLL_R_X71Y126_SLICE_X106Y126_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C3 = CLBLL_L_X2Y124_SLICE_X1Y124_BQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C5 = CLBLL_L_X2Y124_SLICE_X1Y124_DO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_C6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D2 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D3 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D2 = CLBLL_L_X2Y124_SLICE_X1Y124_CQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D3 = CLBLL_L_X2Y124_SLICE_X1Y124_BQ;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D5 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_D6 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_A2 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_L_X2Y124_SLICE_X1Y124_DX = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_A3 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_A4 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_A5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_A6 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_B1 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_B2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_B3 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_B4 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_B5 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_C2 = CLBLM_L_X74Y129_SLICE_X112Y129_F7AMUX_O;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_C3 = CLBLL_R_X73Y129_SLICE_X111Y129_F8MUX_O;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_C4 = CLBLL_R_X73Y129_SLICE_X110Y129_F7AMUX_O;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_C5 = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C5 = LIOB33_X0Y153_IOB_X0Y154_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_C6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_D1 = 1'b1;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_D2 = 1'b1;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_D3 = 1'b1;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_D4 = 1'b1;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_D5 = 1'b1;
  assign CLBLL_R_X73Y129_SLICE_X110Y129_D6 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D2 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D3 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D4 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D5 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_D6 = 1'b1;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_A1 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_A2 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_A3 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_A5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_B1 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_B2 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_B4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_B5 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_B6 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_C1 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_C2 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_C4 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_C5 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_C6 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_L_X70Y121_SLICE_X104Y121_BO6;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X70Y119_SLICE_X105Y119_CO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_D1 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_D2 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_D4 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_D5 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X73Y129_SLICE_X111Y129_D6 = CLBLM_L_X78Y129_SLICE_X120Y129_AO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A2 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A3 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A4 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_A6 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B1 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B2 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B5 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_A3 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_A4 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C1 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C2 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C4 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C5 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_C6 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_A5 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D1 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D2 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D3 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D4 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y121_SLICE_X106Y121_D6 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A1 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A3 = CLBLM_L_X78Y126_SLICE_X120Y126_AO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A4 = CLBLL_R_X79Y124_SLICE_X122Y124_BO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_A6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B2 = CLBLL_R_X77Y129_SLICE_X118Y129_DO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B3 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_CO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B5 = CLBLL_R_X77Y115_SLICE_X118Y115_AO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_B6 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C1 = CLBLM_L_X78Y120_SLICE_X120Y120_CO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C2 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C4 = CLBLL_R_X77Y122_SLICE_X118Y122_BO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_C6 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_A6 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B1 = 1'b1;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D1 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D2 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D4 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D5 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLL_R_X71Y121_SLICE_X107Y121_D6 = CLBLL_R_X77Y113_SLICE_X118Y113_BO6;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B3 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_C3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_B6 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C1 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_C4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C5 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X121Y117_C5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_C6 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X121Y120_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A5 = RIOB33_X105Y57_IOB_X1Y57_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_A6 = LIOB33_X0Y163_IOB_X0Y163_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B3 = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_B6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C1 = LIOB33_X0Y163_IOB_X0Y164_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C2 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C4 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C5 = RIOB33_X105Y57_IOB_X1Y58_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_C6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D1 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D2 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D3 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D4 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D5 = 1'b1;
  assign CLBLM_L_X78Y120_SLICE_X120Y120_D6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_L_X70Y127_SLICE_X104Y127_AO6;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X70Y121_SLICE_X104Y121_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_A1 = CLBLL_R_X71Y121_SLICE_X107Y121_F8MUX_O;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_A2 = CLBLL_R_X71Y121_SLICE_X106Y121_F7AMUX_O;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_A3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_A4 = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_A5 = CLBLL_R_X71Y121_SLICE_X106Y121_F7BMUX_O;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_A6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_B1 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_B2 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_B3 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_B4 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_B5 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_B6 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_B6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_C1 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_C2 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_C3 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_C4 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_C5 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_C6 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_D1 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_D2 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_D3 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_D4 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_D5 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X106Y122_D6 = 1'b1;
  assign CLBLL_R_X75Y119_SLICE_X114Y119_C1 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_C3 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_C4 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_C5 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_A1 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_A2 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_A3 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_A4 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_A5 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_A6 = 1'b1;
  assign CLBLM_L_X78Y117_SLICE_X120Y117_C6 = 1'b1;
  assign CLBLM_L_X72Y125_SLICE_X109Y125_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_B1 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_B2 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_B3 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_B4 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_B5 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_B6 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_C1 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_C2 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_C3 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_C4 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_C5 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_C6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_A6 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_D1 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_D2 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_D3 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_D4 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_D5 = 1'b1;
  assign CLBLL_R_X71Y122_SLICE_X107Y122_D6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_B6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C6 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_C5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D2 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_A6 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X121Y121_D6 = 1'b1;
  assign LIOI3_X0Y203_ILOGIC_X0Y203_D = LIOB33_X0Y203_IOB_X0Y203_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A3 = LIOB33_X0Y165_IOB_X0Y165_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A4 = RIOB33_X105Y59_IOB_X1Y59_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B3 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B1 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_B6 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y80_D = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B2 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C1 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C2 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B3 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_C6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B5 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_L_X70Y123_SLICE_X105Y123_DO6;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D1 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_B6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D2 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D3 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D4 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D5 = 1'b1;
  assign CLBLM_L_X78Y121_SLICE_X120Y121_D6 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign RIOI3_X105Y65_ILOGIC_X1Y66_D = RIOB33_X105Y65_IOB_X1Y66_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y194_D = LIOB33_X0Y193_IOB_X0Y194_I;
  assign LIOI3_TBYTESRC_X0Y193_ILOGIC_X0Y193_D = LIOB33_X0Y193_IOB_X0Y193_I;
  assign RIOI3_X105Y65_ILOGIC_X1Y65_D = RIOB33_X105Y65_IOB_X1Y65_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C1 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C2 = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D3 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C3 = CLBLL_R_X73Y128_SLICE_X110Y128_F8MUX_O;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C4 = CLBLM_L_X72Y128_SLICE_X109Y128_F7AMUX_O;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_C6 = CLBLL_R_X73Y128_SLICE_X111Y128_F7AMUX_O;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D4 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D1 = CLBLM_L_X72Y129_SLICE_X109Y129_F7BMUX_O;
  assign CLBLM_L_X74Y128_SLICE_X113Y128_D6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D4 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D5 = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign CLBLM_L_X72Y128_SLICE_X109Y128_D6 = CLBLL_R_X73Y128_SLICE_X111Y128_F7BMUX_O;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y123_SLICE_X109Y123_C4 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B1 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B2 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A1 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A2 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A3 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A4 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A5 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_A6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B1 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B2 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B3 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B5 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B4 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B5 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_B6 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_B6 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C1 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C2 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C3 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C4 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C5 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_C6 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D1 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D2 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D3 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D4 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D5 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X121Y122_D6 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_D1 = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A3 = RIOB33_X105Y87_IOB_X1Y87_I;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A4 = LIOB33_X0Y193_IOB_X0Y193_I;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A5 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C2 = CLBLL_R_X71Y131_SLICE_X106Y131_CO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_A6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_L_X70Y127_SLICE_X104Y127_BO6;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C3 = CLBLM_L_X72Y129_SLICE_X108Y129_F8MUX_O;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B2 = RIOB33_X105Y59_IOB_X1Y60_I;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_A4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B3 = LIOB33_X0Y165_IOB_X0Y166_I;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C4 = CLBLM_L_X72Y128_SLICE_X108Y128_F7AMUX_O;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B5 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_B6 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C5 = CLBLM_L_X72Y129_SLICE_X109Y129_F7AMUX_O;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C1 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C2 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C3 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C4 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C5 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_C6 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D1 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D2 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D3 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D4 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D5 = 1'b1;
  assign CLBLM_L_X78Y122_SLICE_X120Y122_D6 = 1'b1;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_B1 = CLBLM_L_X70Y121_SLICE_X104Y121_DQ;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D1 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D2 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D3 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D4 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D5 = 1'b1;
  assign CLBLM_L_X72Y128_SLICE_X108Y128_D6 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C4 = 1'b1;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A5 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_C6 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_B6 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y167_ILOGIC_X1Y168_D = RIOB33_X105Y167_IOB_X1Y168_I;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D1 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C4 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D2 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X70Y123_SLICE_X104Y123_D3 = 1'b1;
  assign CLBLM_L_X74Y123_SLICE_X113Y123_C6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign RIOI3_X105Y71_ILOGIC_X1Y72_D = RIOB33_X105Y71_IOB_X1Y72_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y71_ILOGIC_X1Y71_D = RIOB33_X105Y71_IOB_X1Y71_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLM_L_X74Y128_SLICE_X112Y128_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A1 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A2 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A3 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A4 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A5 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_A6 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B1 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B2 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B3 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B4 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B5 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_B6 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C1 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C2 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C3 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C4 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C5 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_C6 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_L_X70Y127_SLICE_X104Y127_DO6;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C3 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D1 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D2 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D3 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D4 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D5 = 1'b1;
  assign CLBLM_L_X78Y123_SLICE_X121Y123_D6 = 1'b1;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_C6 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A2 = RIOB33_X105Y189_IOB_X1Y190_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A5 = RIOB33_X105Y73_IOB_X1Y74_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_A6 = LIOB33_X0Y179_IOB_X0Y180_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B5 = RIOB33_X105Y85_IOB_X1Y86_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_B6 = LIOB33_X0Y191_IOB_X0Y192_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C2 = LIOB33_SING_X0Y199_IOB_X0Y199_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C4 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_C6 = RIOB33_X105Y93_IOB_X1Y93_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D1 = LIOB33_X0Y171_IOB_X0Y171_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D2 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D5 = RIOB33_X105Y65_IOB_X1Y65_I;
  assign CLBLM_L_X78Y123_SLICE_X120Y123_D6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X72Y118_SLICE_X109Y118_D1 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B4 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_B6 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C4 = CLBLM_L_X74Y125_SLICE_X112Y125_F7AMUX_O;
  assign RIOI3_X105Y189_ILOGIC_X1Y190_D = RIOB33_X105Y189_IOB_X1Y190_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y84_D = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A5 = CLBLM_L_X78Y123_SLICE_X120Y123_BO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOI3_X0Y83_ILOGIC_X0Y83_D = LIOB33_X0Y83_IOB_X0Y83_I;
  assign RIOI3_X105Y189_ILOGIC_X1Y189_D = RIOB33_X105Y189_IOB_X1Y189_I;
  assign CLBLM_L_X72Y118_SLICE_X108Y118_A6 = CLBLL_R_X73Y119_SLICE_X111Y119_DO6;
  assign CLBLM_L_X74Y123_SLICE_X112Y123_C6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A1 = CLBLL_R_X71Y126_SLICE_X107Y126_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A2 = CLBLL_R_X71Y125_SLICE_X107Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A3 = CLBLL_R_X71Y127_SLICE_X107Y127_AO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A4 = CLBLL_R_X75Y125_SLICE_X115Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A5 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_A6 = CLBLM_L_X72Y128_SLICE_X108Y128_CO6;
  assign RIOI3_X105Y67_ILOGIC_X1Y68_D = RIOB33_X105Y67_IOB_X1Y68_I;
  assign RIOI3_X105Y67_ILOGIC_X1Y67_D = RIOB33_X105Y67_IOB_X1Y67_I;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B1 = CLBLL_R_X71Y126_SLICE_X107Y126_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B2 = CLBLL_R_X71Y125_SLICE_X107Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B3 = CLBLL_R_X71Y127_SLICE_X107Y127_AO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B4 = CLBLL_R_X75Y125_SLICE_X115Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B5 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_B6 = CLBLM_L_X72Y128_SLICE_X108Y128_CO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C1 = CLBLL_R_X71Y127_SLICE_X107Y127_AO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C2 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C3 = CLBLL_R_X71Y125_SLICE_X107Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C4 = CLBLM_L_X72Y128_SLICE_X108Y128_CO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C5 = CLBLL_R_X71Y126_SLICE_X107Y126_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_C6 = CLBLL_R_X75Y125_SLICE_X115Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D1 = CLBLL_R_X71Y127_SLICE_X107Y127_AO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D2 = CLBLL_R_X71Y125_SLICE_X107Y125_CO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D3 = CLBLL_R_X71Y125_SLICE_X107Y125_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D4 = CLBLM_L_X72Y128_SLICE_X108Y128_CO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D5 = CLBLL_R_X71Y126_SLICE_X107Y126_DO6;
  assign CLBLL_R_X71Y125_SLICE_X106Y125_D6 = CLBLL_R_X75Y125_SLICE_X115Y125_DO6;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A1 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A5 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_A6 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B1 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B3 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B5 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_B6 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C1 = CLBLM_L_X56Y116_SLICE_X84Y116_CO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C3 = CLBLL_R_X73Y125_SLICE_X110Y125_F8MUX_O;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C4 = CLBLL_R_X71Y125_SLICE_X107Y125_F7AMUX_O;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C5 = CLBLM_L_X72Y125_SLICE_X108Y125_F7AMUX_O;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_C6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D1 = CLBLM_L_X72Y125_SLICE_X108Y125_F7BMUX_O;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D4 = CLBLM_L_X72Y125_SLICE_X109Y125_F8MUX_O;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D5 = CLBLM_L_X72Y124_SLICE_X108Y124_F7AMUX_O;
  assign CLBLL_R_X71Y125_SLICE_X107Y125_D6 = CLBLM_L_X70Y128_SLICE_X104Y128_BO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_A6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_B6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_C6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X121Y124_D6 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A4 = LIOB33_X0Y185_IOB_X0Y185_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A5 = RIOB33_X105Y79_IOB_X1Y79_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_A6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B2 = RIOB33_X105Y81_IOB_X1Y82_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B5 = LIOB33_X0Y187_IOB_X0Y188_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_B6 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_C6 = 1'b1;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D1 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D2 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D3 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D4 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D5 = 1'b1;
  assign CLBLM_L_X78Y124_SLICE_X120Y124_D6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X74Y126_SLICE_X112Y126_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_A1 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_A2 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_A3 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_A4 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_A5 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_A6 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_B1 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_B2 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_B3 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_B4 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_B5 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_B6 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_C1 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_C2 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_C3 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_C4 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_C5 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_C6 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_D1 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_D2 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_D3 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_D4 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_D5 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X85Y116_D6 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_A1 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_A3 = CLBLM_L_X56Y116_SLICE_X84Y116_AQ;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_A4 = CLBLM_L_X56Y116_SLICE_X84Y116_BO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_A5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_A6 = CLBLL_R_X71Y116_SLICE_X107Y116_BO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_AX = CLBLM_L_X56Y116_SLICE_X84Y116_CO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_B2 = CLBLM_L_X56Y116_SLICE_X84Y116_BQ;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_B3 = CLBLM_L_X56Y116_SLICE_X84Y116_AQ;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_B6 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_BX = CLBLM_L_X56Y116_SLICE_X84Y116_AO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_C1 = CLBLM_L_X56Y116_SLICE_X84Y116_BQ;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_C2 = CLBLM_L_X56Y116_SLICE_X84Y116_AQ;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_C3 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_C5 = RIOB33_X105Y165_IOB_X1Y165_I;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_C6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A1 = CLBLL_R_X75Y125_SLICE_X115Y125_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A2 = CLBLL_R_X75Y125_SLICE_X114Y125_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A3 = CLBLL_R_X71Y126_SLICE_X107Y126_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A4 = CLBLL_R_X73Y127_SLICE_X111Y127_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A5 = CLBLM_L_X74Y125_SLICE_X112Y125_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_A6 = CLBLM_L_X72Y124_SLICE_X108Y124_CO6;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_D3 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_D1 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_D6 = 1'b1;
  assign CLBLM_L_X56Y116_SLICE_X84Y116_D2 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B1 = CLBLL_R_X75Y125_SLICE_X115Y125_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B2 = CLBLL_R_X75Y125_SLICE_X114Y125_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B3 = CLBLL_R_X71Y126_SLICE_X107Y126_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B4 = CLBLM_L_X72Y124_SLICE_X108Y124_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B5 = CLBLM_L_X74Y125_SLICE_X112Y125_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_B6 = CLBLL_R_X73Y127_SLICE_X111Y127_CO6;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C1 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C2 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C3 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C4 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C5 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_C6 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D1 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D2 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D3 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D4 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D5 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X106Y126_D6 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A1 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A2 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A3 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_A6 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B1 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_CO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B4 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_B6 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLL_L_X2Y124_SLICE_X1Y124_AO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C1 = CLBLL_R_X73Y126_SLICE_X111Y126_F7BMUX_O;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C2 = CLBLM_L_X72Y126_SLICE_X109Y126_F7AMUX_O;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C3 = CLBLL_R_X73Y126_SLICE_X110Y126_F8MUX_O;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C4 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_C6 = CLBLM_L_X70Y124_SLICE_X105Y124_BO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D1 = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D2 = CLBLM_L_X72Y126_SLICE_X108Y126_F8MUX_O;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D3 = CLBLM_L_X72Y126_SLICE_X109Y126_F7BMUX_O;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D4 = CLBLL_R_X71Y126_SLICE_X107Y126_F7AMUX_O;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X71Y126_SLICE_X107Y126_D6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_L_X70Y121_SLICE_X105Y121_CO6;
  assign CLBLM_L_X72Y125_SLICE_X108Y125_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_D1 = CLBLM_L_X70Y119_SLICE_X104Y119_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_L_X2Y123_SLICE_X0Y123_DO6;
  assign LIOI3_X0Y85_OLOGIC_X0Y86_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A1 = CLBLL_R_X73Y127_SLICE_X111Y127_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A2 = CLBLM_L_X72Y124_SLICE_X108Y124_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A3 = CLBLM_L_X74Y125_SLICE_X112Y125_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A4 = CLBLL_R_X75Y125_SLICE_X115Y125_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A5 = CLBLL_R_X75Y125_SLICE_X114Y125_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_A6 = CLBLL_R_X71Y126_SLICE_X107Y126_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B1 = CLBLL_R_X73Y127_SLICE_X111Y127_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B2 = CLBLM_L_X72Y124_SLICE_X108Y124_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B3 = CLBLM_L_X74Y125_SLICE_X112Y125_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B4 = CLBLL_R_X75Y125_SLICE_X115Y125_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B5 = CLBLL_R_X75Y125_SLICE_X114Y125_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_B6 = CLBLL_R_X71Y126_SLICE_X107Y126_CO6;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_C6 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X106Y127_D6 = 1'b1;
  assign RIOI3_X105Y95_ILOGIC_X1Y96_D = RIOB33_X105Y95_IOB_X1Y96_I;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLL_L_X2Y124_SLICE_X0Y124_AO6;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X2Y123_SLICE_X1Y123_AO6;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A1 = CLBLM_L_X72Y127_SLICE_X109Y127_F8MUX_O;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A2 = CLBLM_L_X72Y127_SLICE_X108Y127_F7AMUX_O;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A4 = CLBLM_L_X72Y127_SLICE_X108Y127_F7BMUX_O;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A5 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_A6 = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign RIOI3_X105Y95_ILOGIC_X1Y95_D = RIOB33_X105Y95_IOB_X1Y95_I;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_B6 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_C6 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_D4 = 1'b1;
  assign RIOI3_X105Y191_ILOGIC_X1Y192_D = RIOB33_X105Y191_IOB_X1Y192_I;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_D5 = 1'b1;
  assign RIOI3_X105Y191_ILOGIC_X1Y191_D = RIOB33_X105Y191_IOB_X1Y191_I;
  assign LIOI3_X0Y85_ILOGIC_X0Y85_D = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_D6 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D1 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D2 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D3 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D4 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D5 = 1'b1;
  assign CLBLL_R_X71Y127_SLICE_X107Y127_D6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_A2 = RIOB33_X105Y61_IOB_X1Y61_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_A3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_A4 = LIOB33_X0Y167_IOB_X0Y167_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_A5 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_A6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_A1 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_A2 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_B2 = LIOB33_X0Y185_IOB_X0Y186_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_B3 = RIOB33_X105Y79_IOB_X1Y80_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_B5 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_B6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_A3 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_A4 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_A5 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_C1 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_C2 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_C3 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_C4 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_C5 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_C6 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_B2 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_B3 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_B4 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_B5 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_B6 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_C1 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_C2 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_D1 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_D2 = 1'b1;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_A6 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_D3 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_D4 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_D5 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X122Y123_D6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A4 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_D1 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A5 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_D2 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_D3 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_D4 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_D5 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_A6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X78Y126_SLICE_X121Y126_D6 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_A1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_A3 = LIOB33_X0Y187_IOB_X0Y187_I;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_A4 = RIOB33_X105Y81_IOB_X1Y81_I;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_A5 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C3 = CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_A6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C4 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_B1 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_B2 = LIOB33_X0Y181_IOB_X0Y181_I;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B2 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C5 = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_A1 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_A2 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_A3 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_A4 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_A5 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_A6 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_B3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B4 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_B1 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_B2 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_B3 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_B4 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_B5 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_B6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_B6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B3 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_C1 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_C2 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_C3 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_C4 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_C5 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_C6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B4 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B5 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_D1 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_D2 = 1'b1;
  assign CLBLM_L_X78Y126_SLICE_X120Y126_D3 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_B6 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_D1 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_D2 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_D3 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_D4 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_D5 = 1'b1;
  assign CLBLL_R_X79Y123_SLICE_X123Y123_D6 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_B5 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_C1 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_B6 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C2 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C3 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C4 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C5 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_C6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_A1 = CLBLL_R_X77Y129_SLICE_X118Y129_CO6;
  assign CLBLL_R_X77Y122_SLICE_X119Y122_D1 = 1'b1;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_A2 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A1 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A2 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_A3 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A3 = CLBLL_R_X71Y128_SLICE_X106Y128_AQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A4 = CLBLL_R_X71Y128_SLICE_X106Y128_BO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A5 = CLBLL_R_X71Y127_SLICE_X106Y127_BO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_A6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_A4 = CLBLM_L_X78Y123_SLICE_X120Y123_AO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_AX = CLBLL_R_X71Y128_SLICE_X106Y128_CO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D1 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B1 = RIOB33_X105Y153_IOB_X1Y154_I;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B2 = CLBLL_R_X71Y128_SLICE_X106Y128_BQ;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_A5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B3 = CLBLL_R_X71Y128_SLICE_X106Y128_AQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_B6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_A6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_BX = CLBLL_R_X71Y128_SLICE_X106Y128_AO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D2 = CLBLM_L_X78Y120_SLICE_X120Y120_AO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C1 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C2 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C3 = CLBLL_R_X71Y128_SLICE_X106Y128_AQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C4 = RIOB33_X105Y155_IOB_X1Y155_I;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C5 = CLBLL_R_X71Y128_SLICE_X106Y128_BQ;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_C6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D3 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D4 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X2Y124_SLICE_X0Y124_CO6;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X2Y124_SLICE_X1Y124_CO6;
  assign CLBLM_L_X72Y129_SLICE_X109Y129_D6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X106Y128_D6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_B1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_B2 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_B3 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_B4 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_B5 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLL_R_X75Y120_SLICE_X115Y120_B6 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_A6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A1 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_B6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D1 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_C6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A5 = CLBLM_L_X78Y119_SLICE_X120Y119_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_A6 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLL_R_X77Y131_SLICE_X119Y131_C4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D1 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D2 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D3 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D4 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D5 = 1'b1;
  assign CLBLL_R_X71Y128_SLICE_X107Y128_D6 = 1'b1;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D2 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_A2 = RIOB33_X105Y61_IOB_X1Y62_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_A3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_A4 = LIOB33_X0Y167_IOB_X0Y168_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_A5 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_A6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_B5 = CLBLL_R_X73Y119_SLICE_X111Y119_CO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_B2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_B3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_B4 = RIOB33_X105Y67_IOB_X1Y67_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_B5 = LIOB33_X0Y173_IOB_X0Y173_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_B6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_B6 = CLBLM_L_X70Y117_SLICE_X105Y117_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B1 = CLBLM_L_X76Y131_SLICE_X116Y131_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B2 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_C1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_C2 = RIOB33_X105Y65_IOB_X1Y66_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_C3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_C4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_C5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_C6 = LIOB33_X0Y171_IOB_X0Y172_I;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D3 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B3 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B4 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B5 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_D1 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_D2 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_D3 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_D4 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_D5 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X122Y124_D6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y123_SLICE_X108Y123_D4 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_C5 = CLBLM_L_X72Y118_SLICE_X108Y118_DO6;
  assign RIOI3_X105Y155_ILOGIC_X1Y156_D = RIOB33_X105Y155_IOB_X1Y156_I;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X68Y119_SLICE_X103Y119_C6 = CLBLM_L_X72Y118_SLICE_X108Y118_CO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C1 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_A1 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_A2 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_A3 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_A4 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_A5 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_A6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C2 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign RIOI3_X105Y155_ILOGIC_X1Y155_D = RIOB33_X105Y155_IOB_X1Y155_I;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_B1 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_B2 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_B3 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_B4 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_B5 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_B6 = 1'b1;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C4 = CLBLM_L_X78Y117_SLICE_X120Y117_BO6;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_C1 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_C2 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_C3 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_C4 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_C5 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_C6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_A6 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C5 = CLBLM_L_X98Y132_SLICE_X154Y132_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_C6 = CLBLM_L_X76Y131_SLICE_X116Y131_BO6;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_D1 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_D2 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_D3 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_D4 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_D5 = 1'b1;
  assign CLBLL_R_X79Y124_SLICE_X123Y124_D6 = 1'b1;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B1 = RIOB33_X105Y159_IOB_X1Y160_I;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B2 = CLBLM_L_X70Y124_SLICE_X104Y124_BQ;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B3 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X70Y124_SLICE_X104Y124_B4 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D1 = CLBLL_R_X77Y130_SLICE_X118Y130_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D2 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D3 = CLBLL_R_X77Y130_SLICE_X118Y130_BO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign CLBLM_L_X72Y129_SLICE_X108Y129_D6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A1 = CLBLL_R_X73Y129_SLICE_X110Y129_CO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A2 = CLBLL_R_X75Y127_SLICE_X114Y127_CO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A3 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A4 = CLBLM_L_X74Y128_SLICE_X112Y128_CO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A5 = CLBLM_L_X72Y128_SLICE_X109Y128_DO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_A6 = CLBLM_L_X72Y128_SLICE_X109Y128_CO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X2Y124_SLICE_X0Y124_DO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B2 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B3 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B5 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_B6 = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_D1 = CLBLL_R_X71Y128_SLICE_X106Y128_AO6;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C2 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C3 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C5 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_C6 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_B6 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign LIOI3_X0Y89_OLOGIC_X0Y90_T1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D2 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D3 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D5 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X106Y129_D6 = 1'b1;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_D1 = CLBLM_L_X70Y128_SLICE_X105Y128_CO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_C1 = CLBLM_L_X78Y117_SLICE_X120Y117_AO6;
  assign LIOI3_X0Y89_OLOGIC_X0Y89_T1 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_C2 = CLBLL_R_X77Y113_SLICE_X118Y113_AO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_C3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A2 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A3 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A5 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_A6 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_C5 = CLBLL_R_X77Y129_SLICE_X118Y129_AO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_C6 = CLBLL_R_X79Y125_SLICE_X122Y125_AO6;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B2 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B3 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B5 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_B6 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C2 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C3 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C5 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_C6 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D1 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D2 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D3 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D4 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D5 = 1'b1;
  assign CLBLL_R_X71Y129_SLICE_X107Y129_D6 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_A2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_A3 = LIOB33_X0Y169_IOB_X0Y170_I;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_A4 = RIOB33_X105Y63_IOB_X1Y64_I;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_A5 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_A6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_B1 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_B2 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_B3 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_B4 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_B5 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_B6 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_D1 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_D2 = CLBLL_R_X77Y130_SLICE_X118Y130_CO6;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_C1 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_C2 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_C3 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_C4 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_C5 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_C6 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_D3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_D4 = CLBLM_L_X78Y120_SLICE_X120Y120_BO6;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_D5 = CLBLL_R_X79Y123_SLICE_X122Y123_AO6;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_D1 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_D2 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_D3 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_D4 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_D5 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X122Y125_D6 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X113Y124_D6 = CLBLL_R_X77Y131_SLICE_X118Y131_BO6;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_A1 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_A2 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_A3 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_A4 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_A5 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_A6 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_A1 = CLBLL_R_X77Y131_SLICE_X118Y131_DO6;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_B1 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_B2 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_B3 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_B4 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_B5 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_B6 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_A3 = CLBLL_R_X77Y131_SLICE_X118Y131_AO6;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_C1 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_C2 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_C3 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_C4 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_C5 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_C6 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_A4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_A5 = CLBLM_L_X76Y133_SLICE_X117Y133_AO6;
  assign LIOI3_X0Y151_ILOGIC_X0Y152_D = LIOB33_X0Y151_IOB_X0Y152_I;
  assign LIOI3_X0Y151_ILOGIC_X0Y151_D = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_A6 = CLBLM_L_X78Y119_SLICE_X120Y119_CO6;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_D1 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_D2 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_D3 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_D4 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_D5 = 1'b1;
  assign CLBLL_R_X79Y125_SLICE_X123Y125_D6 = 1'b1;
  assign RIOI3_X105Y195_ILOGIC_X1Y196_D = RIOB33_X105Y195_IOB_X1Y196_I;
  assign RIOI3_X105Y195_ILOGIC_X1Y195_D = RIOB33_X105Y195_IOB_X1Y195_I;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_B1 = CLBLM_L_X98Y131_SLICE_X154Y131_AO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_B2 = CLBLL_R_X79Y124_SLICE_X122Y124_AO6;
  assign RIOI3_X105Y73_ILOGIC_X1Y74_D = RIOB33_X105Y73_IOB_X1Y74_I;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_D1 = CLBLL_R_X71Y131_SLICE_X106Y131_CO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_B3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign RIOI3_X105Y73_ILOGIC_X1Y73_D = RIOB33_X105Y73_IOB_X1Y73_I;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_B4 = CLBLL_R_X77Y133_SLICE_X118Y133_BO6;
  assign LIOI3_SING_X0Y99_OLOGIC_X0Y99_T1 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_B5 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_B6 = CLBLM_L_X78Y119_SLICE_X120Y119_BO6;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X2Y123_SLICE_X0Y123_CO6;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y158_D = RIOB33_X105Y157_IOB_X1Y158_I;
  assign RIOI3_TBYTESRC_X105Y157_ILOGIC_X1Y157_D = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_C2 = CLBLL_R_X77Y133_SLICE_X118Y133_AO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_C4 = CLBLM_L_X76Y127_SLICE_X116Y127_CO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_C5 = CLBLL_R_X77Y130_SLICE_X118Y130_DO6;
  assign CLBLM_L_X74Y124_SLICE_X112Y124_C6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_B4 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_B5 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_B6 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_C1 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_C2 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_C3 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_C4 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_C5 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_C6 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_C3 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X2Y123_SLICE_X0Y123_AO6;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A1 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_C4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A5 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_C5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_A6 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_D1 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_C6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_B6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_C6 = 1'b1;
  assign CLBLL_R_X77Y133_SLICE_X119Y133_D6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X121Y129_D6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A3 = LIOB33_X0Y173_IOB_X0Y174_I;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A5 = RIOB33_X105Y67_IOB_X1Y68_I;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_A6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B1 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_D1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B5 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_D2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_B6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C1 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_D3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C5 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_D4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_C6 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_D5 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D2 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X117Y131_D6 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D1 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D2 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D3 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D4 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D5 = 1'b1;
  assign CLBLM_L_X78Y129_SLICE_X120Y129_D6 = 1'b1;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D3 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_A1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_A2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D4 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_A3 = LIOB33_X0Y183_IOB_X0Y184_I;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_A4 = RIOB33_X105Y77_IOB_X1Y78_I;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_A6 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D5 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLM_R_X59Y118_SLICE_X88Y118_AO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A1 = CLBLL_R_X71Y131_SLICE_X106Y131_DO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A2 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A3 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A4 = CLBLL_R_X71Y131_SLICE_X106Y131_BO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A5 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_A6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_AX = CLBLL_R_X71Y131_SLICE_X106Y131_CO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_B1 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B1 = CLBLL_R_X71Y131_SLICE_X106Y131_BQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B2 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B3 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B4 = RIOB33_X105Y161_IOB_X1Y162_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B5 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_B6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_B2 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X76Y133_SLICE_X117Y133_D6 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_BX = CLBLL_R_X71Y131_SLICE_X106Y131_AO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_B3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C1 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C2 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C3 = CLBLL_R_X71Y131_SLICE_X106Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C4 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C5 = CLBLL_R_X71Y131_SLICE_X106Y131_BQ;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_C6 = RIOB33_X105Y163_IOB_X1Y163_I;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_B4 = LIOB33_X0Y197_IOB_X0Y198_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_B5 = RIOB33_X105Y91_IOB_X1Y92_I;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_B6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D1 = CLBLM_L_X72Y128_SLICE_X109Y128_DO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D2 = CLBLL_R_X75Y128_SLICE_X115Y128_CO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D3 = CLBLL_R_X73Y129_SLICE_X110Y129_CO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D4 = CLBLM_L_X74Y128_SLICE_X112Y128_CO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D5 = CLBLL_R_X75Y127_SLICE_X114Y127_CO6;
  assign CLBLL_R_X71Y131_SLICE_X106Y131_D6 = CLBLM_L_X72Y128_SLICE_X109Y128_CO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_C1 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_C2 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A1 = RIOB33_X105Y171_IOB_X1Y171_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A2 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A3 = CLBLL_R_X71Y131_SLICE_X107Y131_CQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A4 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A5 = CLBLM_L_X72Y131_SLICE_X108Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_A6 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_C3 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_AX = CLBLL_R_X71Y131_SLICE_X107Y131_DO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B1 = CLBLL_R_X71Y131_SLICE_X107Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B2 = CLBLM_L_X72Y131_SLICE_X108Y131_CO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B3 = LIOB33_X0Y81_IOB_X0Y82_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B4 = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B5 = CLBLL_R_X71Y131_SLICE_X107Y131_CO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_B6 = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_C4 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_C5 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C3 = RIOB33_X105Y155_IOB_X1Y156_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C4 = CLBLL_R_X71Y131_SLICE_X107Y131_BQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C5 = CLBLL_R_X71Y131_SLICE_X107Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_C6 = CLBLM_L_X44Y118_SLICE_X66Y118_AO6;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_C6 = 1'b1;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X1Y32_O;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_CX = CLBLM_L_X72Y131_SLICE_X108Y131_AO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D1 = CLBLM_L_X46Y116_SLICE_X70Y116_AO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D2 = CLBLM_L_X46Y116_SLICE_X70Y116_BO6;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D3 = RIOB33_X105Y157_IOB_X1Y157_I;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D4 = CLBLL_R_X71Y131_SLICE_X107Y131_BQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D5 = CLBLL_R_X71Y131_SLICE_X107Y131_AQ;
  assign CLBLL_R_X71Y131_SLICE_X107Y131_D6 = CLBLM_R_X49Y116_SLICE_X74Y116_AO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B2 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B3 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B4 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_D1 = CLBLL_R_X71Y131_SLICE_X107Y131_BO6;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B5 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_D1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_B6 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_D2 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y92_T1 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_D3 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_D4 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_A1 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_A2 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_A3 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_A4 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_A5 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_A6 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_D5 = 1'b1;
  assign CLBLM_L_X76Y131_SLICE_X116Y131_D6 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_B1 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_B2 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_B3 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_B4 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_B5 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_B6 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C2 = 1'b1;
  assign LIOI3_X0Y91_OLOGIC_X0Y91_T1 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_C1 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_C2 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_C3 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_C4 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_C5 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_C6 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C3 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C4 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_C5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A3 = LIOB33_X0Y155_IOB_X0Y156_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A5 = RIOB33_SING_X105Y50_IOB_X1Y50_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_A6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_D1 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_D2 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X117Y120_D3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_B6 = LIOB33_X0Y151_IOB_X0Y151_I;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_A1 = CLBLL_R_X77Y122_SLICE_X118Y122_CO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_A2 = CLBLL_R_X77Y114_SLICE_X118Y114_BO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_A3 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C2 = LIOB33_SING_X0Y150_IOB_X0Y150_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C3 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C4 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_C6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_A4 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_A5 = CLBLL_R_X77Y122_SLICE_X118Y122_AO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_A6 = CLBLM_L_X78Y126_SLICE_X120Y126_BO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_AX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_B1 = CLBLM_L_X78Y124_SLICE_X120Y124_AO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_B2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_B3 = CLBLM_L_X78Y123_SLICE_X120Y123_DO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_B4 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D1 = LIOB33_X0Y151_IOB_X0Y152_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D2 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D3 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_R_X77Y113_SLICE_X118Y113_D6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_BX = LIOB33_X0Y81_IOB_X0Y81_I;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_C1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_C2 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X72Y124_SLICE_X108Y124_D6 = 1'b1;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_C3 = CLBLL_R_X77Y114_SLICE_X118Y114_AO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_C4 = CLBLM_L_X78Y122_SLICE_X120Y122_BO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_C5 = CLBLL_R_X77Y113_SLICE_X118Y113_DO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_C6 = CLBLM_L_X78Y123_SLICE_X120Y123_CO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_CX = LIOB33_X0Y79_IOB_X0Y80_I;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_D1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_D2 = CLBLL_R_X77Y122_SLICE_X118Y122_DO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_D3 = CLBLL_R_X75Y118_SLICE_X114Y118_DO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_D4 = CLBLL_R_X79Y123_SLICE_X122Y123_BO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_D5 = CLBLM_L_X78Y122_SLICE_X120Y122_AO6;
  assign CLBLM_L_X76Y120_SLICE_X116Y120_D6 = CLBLL_R_X79Y124_SLICE_X122Y124_CO6;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_A6 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D5 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X121Y119_D6 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_C6 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D1 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D2 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D3 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D4 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D5 = 1'b1;
  assign CLBLL_R_X77Y113_SLICE_X119Y113_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A2 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A3 = LIOB33_X0Y159_IOB_X0Y160_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y154_D = LIOB33_X0Y153_IOB_X0Y154_I;
  assign LIOI3_X0Y153_ILOGIC_X0Y153_D = LIOB33_X0Y153_IOB_X0Y153_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A5 = RIOB33_X105Y53_IOB_X1Y54_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_A6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign RIOI3_X105Y197_ILOGIC_X1Y198_D = RIOB33_X105Y197_IOB_X1Y198_I;
  assign RIOI3_X105Y197_ILOGIC_X1Y197_D = RIOB33_X105Y197_IOB_X1Y197_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y75_ILOGIC_X1Y76_D = RIOB33_X105Y75_IOB_X1Y76_I;
  assign RIOI3_X105Y75_ILOGIC_X1Y75_D = RIOB33_X105Y75_IOB_X1Y75_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B5 = RIOB33_X105Y55_IOB_X1Y56_I;
  assign CLBLM_L_X78Y119_SLICE_X120Y119_B6 = LIOB33_X0Y161_IOB_X0Y162_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y170_D = RIOB33_X105Y169_IOB_X1Y170_I;
  assign RIOI3_TBYTESRC_X105Y169_ILOGIC_X1Y169_D = RIOB33_X105Y169_IOB_X1Y169_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_A1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_A2 = RIOB33_X105Y51_IOB_X1Y52_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_A3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_A4 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_A5 = LIOB33_X0Y157_IOB_X0Y158_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_A6 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_B1 = LIOB33_X0Y83_IOB_X0Y84_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_B3 = LIOB33_X0Y157_IOB_X0Y157_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_B4 = LIOB33_X0Y85_IOB_X0Y85_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_B5 = RIOB33_X105Y51_IOB_X1Y51_I;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_B6 = LIOB33_X0Y83_IOB_X0Y83_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_C1 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_C2 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_C3 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_C4 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_C5 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_C6 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_D1 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_D2 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_D3 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_D4 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_D5 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X118Y114_D6 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_A1 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_A2 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_A3 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_A4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_A5 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_B1 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_B2 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_B3 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_B4 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_B5 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_B6 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_C1 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_C2 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_C3 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_C4 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_C5 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_C6 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_D1 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_D2 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_D3 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_D4 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_D5 = 1'b1;
  assign CLBLL_R_X77Y114_SLICE_X119Y114_D6 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B1 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B2 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B3 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
endmodule
